//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2025 ICLAB FALL Course
//   Lab08       : Testbench and Pattern
//   Author      : Ying-Yu (Inyi) Wang
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : v1.0
//   Note : PATTERN w/ CG (cg_en = 1)
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################



module PATTERN
`protected
6;HaS?YW[4,SLM/G?bZW)L&d=gce<[=d\0^XEWHV8Ca=-TL)0,1#7)]Ng,V?3[:A
.BLJDC_W,2<e=M;g6)V]Z2PXB1dXbG<XK0>S_IM@FOS3#LZ]^BJO9X<=aI2HBLSa
HS4KP[a>^R;H=WdTPcYM20J]T&3RPF,b3W-:X7L7IUb9CN1gK>9.=cP_MOZ1__3W
]_b4D@dF=SFOEgDE_N3Z.\JSS,Y]?Z.&U<JCG+8_=0PBCb;7RBdMd&8DSGY+e.eb
-W.QTJ]-SaC&MLL^\64LU-(2ZSDB2D/]26d2EK8_BMWc@X;3?MS_.3_S/+X4&?QY
36d=FbN.,+)+NJ:BWQ)JFR>cN:P-SJE2@:WCJg9FCTfB9S)+Z1\3=)??G)JU:B67
>I4g0CD2#g0T1(<3Sfg+&b22Q)>XRH;gWZVT),cUF)DDJ&Ve5HM(I\,;80\@V;:e
Mde>aMfQ7]TW8b^N:;IZd/3)^^KCT\gRaJ(D=W9O.XK6FB6HIS^TTRFT_MU7Q0:&
881/TLCeDV2Sde;_A0Ra..K:_9:665ed@[G3K?3<ZK4/^cBbT5T4e;?cY)YJ/2ZY
f&5N_g\P]B6X?E.9WPU=DKI8:E?.40)?CQB1]](?^7#?ZKKJ076C^5cMW5)+ELV1
=2-CHDf2@&C5DM<<CEFSg6JecdY\(Fe#V70/&?N5H8BfO-;1f9,J@3]D;;9>ASXc
0,PBF/G08EV:U6=fIeW.Uee[/+:f2&g68;eT79RFfDa(LJIK2QN67#fWS-b),GDX
HWT)^3f,7BI:IZV.\8&@),OB;fO\>[Z@=/ENE<g97Sf2_?U><KK^XSW0L4,dJR32
>CS]NIX5F04NgY3T1F:4\8,Dd6T(CEQJ:WREH>FI,],+G.1_K#HM6]1f3K>BbgBH
K5[@e]>IaF-fBaCY?cgAG/V/5D0)D:gXc7@E^:YDPF6>f9\GB1=51Q8DU38;<+:,
FT2_U^WK1NL.-C[aW@NHg#bfEPX4-F[PB)_c6W<=KA)^:O#\GVC;fGS5KcM318^<
@+U^VI8ZOH[\;>^3:Y=3=6.SI38.RDNH)@1>2]&/_e\#C:)47XWR1E<V]+AZA2E/
88Y83U,J0Y;Y7:,&;ZQ6JM@bd;[cL&C\ARNc&BDQW__2/Y[G?ISf[TS<4=>S?#=/
VPN21fB,?9&4-M3^b8V\Q;W._+LS,9?Z5R\_WVR9W6]c,U;:L.WB7\YAY7^[+AZR
DD1CD+gG\9Ea[UA6WFPf5c@YSD3Z(6,L8IXC)++-.D;;.-IG=[#TRL1\Q_NS\[R&
WFbV/X#E+eT,9+88]D;_;(=(D?\WV5BaGD4H:9KGf(O_ACUd[#+;R<a+;;K[;2^W
NC;(\0RG-&;Q:7>]d]Ie0cHQOKbB[4V;WeE];FV:1I/D)1[U#dQWcOd;1,]&:Z1(
[7@RW1P^VAg9/O3H4aKM_\JK3>Z?&-A#6O1S]5H_>,VPIW3C62CP.FeZ<9L[Z)F3
11e\QfQ:7Kc=8W?P06#+fG+4;6Q&]QO9PdR-ZFONS>-JQE&K6F7Fe0S+[J8#X4bY
bf@fB3UZSU3WBG0WVD#1@\GLO,^GNH]g?MR0^/JPC0PCa^K>L7CEcL:E,d>YFP)9
;eM>\IE:6<2a1O#,UEG\b/SSH0BS0E373LDDBb21N7_OWW&eV9;AV<3KBGI]TC;V
K=3]?K530KPPB^fd2\Pa,OQa:aGG_8KOC]]IeU_AA]dg,d0AJM@>g86C<B@VY=@S
(&7@@EZ,^)W,d8DE&X84c[2FVW4>:8YJ5]16F>JZ96-ggcS2G#\0_D\EIc>3M(AI
0b&AFGAg::J)4JORR.4UBM6.egWT[KPPg]XT7ZR=#7^3;)gIT/;AcSER-=IGSC/2
ZP,,]1N0:))8:W0Z)e&P[I<?S>QA^?Y2,OPg\ES\.=MHJ/c:;)1)NKW51#>6]MZ5
HN6@J+^HE&MG2=W:5#FA;J9:;>-0R.>;B3JeZ\+Z_Je&7Y:JXA0A=G9X)Q/V:#:P
)?ZH1Ff:+cT/#[2+OX)N:E;QC8BaWQF^BU\&NWQ[T:^]L4_U)V_SfNI?_d5DWN7N
]Q<dQWQfQ]7RY;^0P;/)Ub0;KA.AM50E-bD:/&>f.dP(e>afR5FV7&SV,E_LWUUY
K@a=M>D.@+d4(S2E(?e>]^@0U9..cYKaf\-_V;a1?5-MP(UJBFg,NW#e&d>La?c+
A:DHbDc_OPe=@ZU@]M@G^e_\SZ(Sa?cFKB=&JdBUg82&8ZP8g3/9.BTN5ed:^D6S
)/Za]L.bX++J/>fefW>XY^D[2)^Xd)fCE]^-&(2YFOZU;d7J&OF<O;225Y(=00Dc
.1_CNa@1@\#^G:VeO),TSHE-TS_&P6IJM6.V:O+H^M6TN;>bGR+@ZC=(d-S<Q.,B
GI:O4@_&1C6R;G2-K(<<)&b\NC4N1-K_e^5QOWKf36QFIb=B4AP1L3;,HU0#K&A?
fa-PaFJ:8cJH?fT,U]M^;Z4>@+JK/D[=@O8_6N9@Og/+g_9g+WA)VPN<(-,L47Xb
P/POQ8B?8S4XQb22Q6NK+II?9#=EBAW6YVGgJFU3>5f[<86X[?@FK7=ZJJ+HB1-)
),QG>NeWf)GdM?J7@M^79H+bSe#<[W?_J957RFCDHFMK>\])34.0OVDAIf-Hc(GJ
+7VKb.S&OC>EAGP&^.dgW,^L6IL7Oc;11YdFf)FMe)Ee[,5f4/JA=dD@3@a(OBW<
gfe4V_eXJ,E0;<&U9dY?\U>]2cM)8<Ba?OWe:D@UYJfB=ZKY#[]DI)Ya7S1+XOCT
B5HcECJP\0RebUe>ZMWK_:^KbXTR00E[.+IeV;<89Z^P[S\&Fd\cA0O2>-V5,)gZ
UNC7QGLR]Rc,L>7@SG<?AM9>f]DW^_3.FA_BE;3S2/]S-D>,=^E8a^_XV8C>X0cQ
:d;N1G^V6W)c=^-Q@811DK9@86=6I1?C,]1+TTSQVHNRU5#(F60O28Q;@Y0.0_G#
K0)82>E)XHGMfL7D_E89@;8_f;V:37LVS:EG^<#LR16LRL[F@NVVZNKD@YC(8_\+
gKQ_XaER)DJ>Nd1/)Y2\]8(U8,a[\HZ6O;D26JCK_+Ug.U-0LfU[c,ENO;@7(ACO
8HMMSMS/Cf7G69/88XRf0A8-VM2E?14]-EHLWX2Z-JVB]NY?0HS3_M>(6H:b1^HX
EYS&3):R+TE]D_2^4ef+8g7W.=V#0X?.3+MGGM5F+E1a-XK+RMC)4+&I^1RM68>;
9a/XS9c5DJ)AH/9THOcW5GVH54(6KK,T&N,4fTb\0@O;/Z4PfbI@b)@[)39L0U>M
/\:IU)7/eM5Z&JT2&Xc-SH>>;a#2U;,(MLbA,d,^6Q^?#H[]]FdU_>E3Q])8cXfb
8[8.5W5NG<JM^1a=UR34/:#Y-,Cb>aX(UN)6ONG<AbbYU&38b6B?@KU7R_a0U0E\
9.LZLDPLAa;(YbW()O/KWE2)/=&KOTXY7I>6]RD<QJCFBSS_M7<K#W3:.1RY+^;O
CfX2#F<1g-(U8SP5#@IZ\/P#7QFM+[?=VM66QXK1NR?>&(B?#[_7;5cSI9WIW7-+
QFBN79X9\-a7dM(FTb&:MS_5A;PbG/88RYd-IECN[GKS^5LC.^;.A]9YA)K9G];L
,.b,-PC7\1FeI@FW8JXO4&SDPFB>)C6HF<&&H.4;54P^Sc6Y6DeN1^>Z04dWB4+7
-\;C3M.g)F_6\]DCBHLO47D5NH-Ee\;g_Q^Od.1/c<)d#:BI;e)M_FV-B9K>13Xf
DIbZ0V6_2AN\3e+e153F5]Z;OBQ0[J;_=I.T^^YZTRH<9.?N&d9AQ/JJGQgR[601
Z&[1DZQMbYe9TA@JYMJe-4&C(<fRCT2#a&IHT8+1UG0G5R=[Z=A_OBVWbU3FVCF,
dWAO[<)_@71:Ce1BQJ1P5+[;:_ZPP6UB)fM+K<c,fARP@OAVC+HA=;H)9\RXLISP
UA&AcQ7GR<31^=(e6dc0URcQ^-F2?K6JKEO>O]gUFD=ZXLY1OT>QO78<adeK6Td+
:e7<CJ^GW^#CYGX:3MS]O^I13ZH6SIZB6W0]+7Pa+_N_S6#,NH9bBL_e)g>RNCKH
GF]4BFD[,g3H;=[D8.8\9THK\)KD/D1baWE6.C8^cM5e(fMb95#9e^T4T6=W+I].
DN&T@2-F2;NMLFO;f7b=X]X\[Te0SNMP[c8g-VX&1=<Nb2GNae],E[S=BF)L[4KP
XNM,:d@R\V,7:@.4bC>X<RS;f#GNFe0HBVe)-#+AL;X7>LI)UfA5.0SXQ9fQ4-^U
G:a7CFcSbed4J&f=6&JS?XZ[:NE8@?5M[\_R[@KHO:b5f#IFJOY&>Fa_8-:>;D<7
1-XC-C=CQ@E6.Q6]QfEUW0L5X0VKG7Z;5&&Z,bP&ZX8OHO\fR(R+03b,3?<4>_:T
_D,\]WN,I])g>WPG0H:4Y0/=Y;7P#G<\U&M=VQ_NM6df0N.5#9:IHA]6J<ICdA,M
OZYB/12=+5e=@JVgVVDGH3c(>B7E\)F.+]8_\XNT9Yg,K)_0I],4<R[fa/_5?;c)
gbge+a?/1R.@P:E7[;Ze<99KV/O@.a2g=d-;(/2f6NZJd\4:V+@>?M&IL8)I82;F
KBWFQQ.b/;F<A.HdIc^AO<gcMCVNT9N>FePg_7Ocb#9A&?BH4[S2=/^GZ+:8#TP(
.+-DFEL;:gfDMc<^85NY94]b28?AL=DQG0SH:9)>d>=c\&=f_3E[+;B6,P?e9]J,
&,&_Fa=<C\&H<b\U3Y3BD[^0\N/XRK7eY?J6^L3CAMK8f>d=EGNDVDf-J,12g/1?
IU7_D2/TJC:)cK4MM^.Y5P+NOL(WdJY-7FeT7Ab^<G7<I)4V707Z>X5/?L(<)L:\
#^OaE9NWXKZRA__WBI;F[]O:=_cMZ:Z\8:V5BdO^IaI&G7cPN7E3TP\B()&D4(88
b.0HF&T]1LfQA73;Q&3;^@A>@gb(NQ]H30(4Q]JY)F]B]LNFH@(@BKMD1#=Q@HDT
TZ=F)?YbRcN75Va,7>S#_,+[2Td1XW0:,UPMX[J2)1;)/beF9Y44\>53@9QRTE0J
KAGC)1Q-JQ41H2C#WSZ^;W.PJ+]fB\72^2:b]W14Rd7#;)[0/R[;^^@Z?^9CH:7H
AOXcbYB9F(I+B?4WH;,VN;<ZKfJJBT=U61Z>g+Iabc3-cC#b)252f:^c9R;<4I.8
:63c/0[Q[4dZ.[U8e]1+M61UL=Re)(V[3U\>BXIHTg=\0-_#CKDDORM8eTAZ\a#6
50;=T=7D#a63dgf09P8OMgC7U@DVR1GVgYPUb6T6IG/fSgCGIe66M;;6M=/SR2a=
^Yf8Q(]AAL_FB,-;OTEV4D/Q2]dUIRR(MY&@2c86G?TO)efL3E?B>\/.[bEP5PWA
-QK2T>Q:VfXeFaRS2IF3TDY/Bfg0-LKe+NaK&B:KB)#3RU]5g3a4d)2P1O_4R=5^
T9AGB[_J1+0W#QV(305I;)/38H(&/R&Ce)YDGb>D\Q7&9\^D8]I81#dD9.>c:;Z,
8P)V6?\cH6X]TLA,>6.c4A:Ie=eC1UZ#M0,((/0dBQ\P:d[NCEZT@.L2S_[@YK),
2F7>EGdZ]-:WDW6gS57L3Y.C<-C]C45F\>;_RWK8KIcED,3Se6aXO<&gN^)Vf,1@
_,AJ7(7T)JSP)HT<FOLVK&S=YQ/(Y\gO>8-2f3M_3)3/PN\.e2QF4c\?X9\X/EFT
.a@BE&KPI1ZK]OJ5+N[B67O8+WJE-,4(?LGFXQ-a,#b54/BUFW[IG8B_STg;41)[
5<DF_fN0N5FBJZ3eC72^)B_&8+G<VC(_K(A2>XUdK24=^I\AVE0GQdM>WDdg;+65
1]c;)FE@H-ISX+Y#d<ReCScH4\W\g1Df38:-dAPKT(5e72dQf7P6BF2\ZX)43BZ7
BaS&44aML73M1:UW9#V&ebM6A54c99X[Q6M7#ac2\/DM>UAG+_E<^-KQJ75#T<F2
,GN4R,_,5:#14B^C_::+)CgQfJ0c^eX9B/=II2O/>E&V2,4TWScAeKfVYJ^S4_6N
68#BD/5M0LUJBQ]+Og#2<Fbd?Rb9;f/7V2>>#P^\_7LUddOE/89?\;5@T6Q][2bJ
;d/7CF:H6IMPKJf,HNDHBZ?(GNCce\K@WFf39])b(P>aDFG:_:OU<G4W.9&Z)@\@
.BY2#Y_/^_]Q/^Q(0+N_b9RcN(FF-e-,R^?Y9C3OJE?]NQbNT:C.12Q\VJE:LO]D
C+NHVK,&]F1-&#@gfAefUI8Kd4c6F6]8UGKB-XR8baSL3,O2J2Dd\[dSBWe_[&c8
<.(G?+ca4#998^GYT.R:>3;?MdCVIFFWD0A3IM7_<0XNeVbHQ^2SRVd.<85>0T@)
^;[2L42&P(M+f4FgH1g48V&8bWTU>CagGW8\/4f#43Q<NO4<S0;Ed2=YOOM7ZJ;Q
1&3+dcO)?gG.a>4IbB^B]IG=@5.V#VIC9cAKCbG&@VI-4a,BY[6He9RN:8PRDe<f
QWU(PMK()84AJ8\[SMM^S@8^gC>ET6KZHXC2:LS#ZfQ@0=#D[Z)VNTVOWQ(Bd=;d
_b2a/F\L<0;@:WD]@[PY=8Eb(UI\OfZ[[I_-(d-J=5OC<Y6>._aQ?.RYJReH-Jcf
EZ@A/32M1,HRP^];O?(KN/#Y7G.X;+N3b\7QNg()3NQRXd=I+6(AW-,KS[C]ENge
,_<)e;Q]aX^/Fc5#LH0B^^(L=N0eM&^EZcg.J8^;TGN(#MgYL30U[]&[Q-F06G9Q
:3J5&ffaaX>@&f-cc?4Y7X-a7&LgBDG5<95/HCN0ZXNTHMg,c-c+9=Y0Q7;aQ./,
/WKW[@\GYX/P-JUR>dZgZ#gP^E1420aQBY;NLfZ;^df_K&b8FM=5\:>(&&Y\,G<A
I)WRFRQ7B=g:JS?T^(SF?Y?96FVA0ca8?D0TZ.J9MJ(:8e[ECON4#>7ID,g8agOc
aFA&3GZaV5J>P/bCRbH>I;fBD#?>D0<LQ_1g33D?P3AA,0^K<3Q86/RA_,K[?TV/
B=dC5PeFGR]6<61(IS;Kc0?5MFP=-,=I+CU-Z0/MH=2D/F8FYUKAZ+Va>O[H]LI8
=+K\3aXad;6b0DZK;(4SMDHf:B+PV?QEYG[+B)+I[ZLBQ3aG1OM_SV_V-]W2Y+/Z
[VLX,9_#(6D8(Og?4bfX/B^_UA+6@8?e1P^+9O#VVCIB0<BdU[^DDa^^PWb9Q]c@
S=OR-SMAQ>Y2H#SS>?=,=VeKJRSVN_7,VVZFf6\8T(b-dQ<S+QVb5K<SMJ,\#9]B
6TfZ5FSEgWVa^W@XGC(_CSEdI20+2Y)_>]>DM,]2\KNI2O,g(PCZD(,&CT)OS60g
,FU?;4:-edW:Ad>PP)/JE[@P3..cQ4@;J&>DYKBH(D7bV-\gg?@DL;3SZATX/&WV
L]_SWDGOY)?Pc(-UHH5ec#]PGeEeR#V/6.,b<&T<Z+3eVJHbSXQ-\L^WUGZQ8SN5
KQS5G1a5FD?1]^\2c[MKVZaBTU?Teg,MTMJZ\-7Q8W.Y5d)OH.4)JN)c5.:B:DZ<
2_8GbgY-8,&7,QZ>^aEg7V#])YNR<ZKbG]]17[^TB4O[cb#NNK-S+0,PIHd2RNFC
_=]-,5GJI7\#@9eG1P_M<IX:);ZJPWSb(+E>cIA/V_@gG5(7gNRbO520VX+a<(6&
&d6G7P#X8^:0gTB]GA@D8RV3NA7KPg?HX]UN1RZASe0BK=ZeU,7DGD7</>\OF0W(
Kb?UcXM9^LDR/YZI0\,VOL#AgW&I,-6^;R#37:7A=_E&1:R8f[X#/>K>ecAXL8P^
&e0&NR=@LI;Q/5VbF(RC@040KS1EJL??M^JNFKNIS+;V1(IcA1#HUC:O5-OegB=A
S.TMK4VH(QX=^6KDgRY_RX83R1:#3#BKa,FB;;AF;bZJ&)&fa1.JD;dWAcCS#8?C
DOZfd-&02NLNR6[-W@8M)SWD,1<4X7d@NVc&&g7S>Y]^>=BN8@8g?1X5US_;Q1fa
>#+O@W<;Z4.9FJeLOf&c[dOFdVA(U1DPfJfX+^Y)J-e,HD#-?XW2GWdHgL7?IZf3
f5U<#@L95e@g8/cg,04ScAR0ceVFVBFK1e21d5Z=U:]7<OUYX70Yc8EBL7VV7#JN
+,1>H#<EICUYZX/cb=c+,D>2Nf\/(^@gD>M^b(#H7NI=M[42+4#cLRd/3K8&3CWO
eb>dG8F<54<I4J)(2YFB6_1A<9He7>/S@>29P93BN-)^4Od;1X?d@W@[Ige7:5^f
,#HV9(EJB4M)EP6.:a0W),QV:[&S;>R>;&ORH;32FC13CEG0WZXCDVfdXM\#deT^
S9/\2_6-7bMa)HAOI-3@:,E@)-3f^CQ,E(UU]]\f-]S-Q\T6e;ZH:KaG^F4WV7/4
ZABN7.7YS_bZ?9;S^;&ZCV#\(-[LC&0>F3D1<)>Y[B&Ha#MEI-9]8JN0W4<?-F(A
(d0:?;?;#<:[&bB5S4Od9(K6LB]PcDG9+&U.b)H5\1NdXb;6WdR8#BPHNWg<J)7R
M>?54ZMcRFf&LSAK>F(^aJJ0(ILS312DLWYD4QYe/[;U;Q/Z2,:\:46dN@=16<.?
ZWR:5103+G<11-AIO,0.UJL9BcPEH(;PH-#IHPZMCJXM1>M&Md01U;LM?[UVe&90
G3f/UgW;;X=KT3>DfVLE3Y][1+a<aJ#G;WS#EK)0:QZ?HD/b9I4_<LC_9[2e9ce/
M-^Y,?-A4Q^\LeER]8881O;;22]g[\H#[abAL<L2I^:./IK(a(K9+JVY(Nca89I<
3&FMZ_UR^Z@#AWM1gK)&IW-(_a@.A.,3A#FGDP^/VG35dCAa150aJ==U7)C:9#.4
_FW<f=ecA<f;^\agaaAY/\992<KgZ\GUA>[1)7eDW(Q8cHA#BI-a5VaX@&C\VRX\
X91M1GUdFP_CfONYe06H)4(#JZ\f^J(.eJ=K>4QND&,-U5RgR<gW.Y.-<^W5\G6#
K@K(4K&,;b7bKfZ_)Q[PT,6FB+/H\,ca[^E.a,T0VXDP_Z(Y/X?8D>bBRG,_B4Y=
H:bbHOO7;Qe@+UeB;Z9N.S#HfP&MD0C8+2GNZ@@]U:VE5>L;I,-U7;G0>\S\BU^A
?I2f34?P]QA@V-#VZT<+__G=R\:DT#=dZ]A?>5PIYU,KJWAVd6ZV&c_0N6_X.d8b
DZW-8=82fC#.eS;ZFH)(D9DB[ODD:1UTBLJJYI^^@[SE3^3CAH_Ue:D-U,W[HS.a
4QV?DG#+57Dd[F8)8EK\+QcX-SH/B:2b1AB7[S2-7aG0IU@U1C7e2F<UT1<Gaf5+
#@9S_Z3J,Z=>(B_bAW7Y&A4.5XRQe22gK@E7QSMD(8G:;/8>D:g2ZJ)9TL@A[VZ,
Ua])J/(7/Z<Q,a.^CV)&-<X#[__QfKK5,/YODA,KL<C,T@2A00\),eDYBIKY,MZ+
W=H6Z\fDA[<G0PO-Q6^V^gC,0bIOQ26=SB:U+7?DC[8]^=A[=f06;ZHES/:N/Saa
#Z#a[PaTOg^DDSFA;;_MESONV8JG7[HDF@HE>]9aWF,>6@V>B9DR&B#7^U\)bQHP
gL98eM90F[7TFM2<@RF1FcTK=]1a[5+e1OG7&H@6.NQ&@=8[=]cMSF&T3#W87SYO
(+fPc_JA/SKV#7-.[\07MJLER6LE<UWHD^6E5/?7\&6&&<TKYZ@R38(1LZUgLO-O
04#I0EWQ-2#4I_..+0(1NMa-5NUf2WKJ(#SVHI_<V:<bNa+bOZY[cc[B]25R>5bG
KVG#OW;WS4JaWY-0+@/_2J8.7:fD&-C,IH\e86XMLVJPP+BbR2.^3&aA8f^W]X0>
U1P5034aBM[[YA8<8A+4F,WIOZAWMbW6d?L\>5]+RIT+1KQ/F<Z:GX6X>a>YdG:X
+K((H0PaVB/g>[2[4\0W55-I]9C:7.M[T9V/b81f\/1+a=FOUUeZ//EWUP@6WQ<f
fE^L5^\>_6(459_K64;SC^<D>5Q-T9F,0,(^,#GRHMcS\cKQb8._^HC\>GR;Q1=4
9/d6a_3b@:?KN1WEfE8bIB7aaHU,C3N4#W,GKgcg7)[cLWc[14IU@W+2eW1)+J&g
EQMg3H]8e98QJT5B=U710,5O]b1=VB5,LXf,3c&TVIYSC2HWH6H.3c^]-Wd^:,>6
QBZ:0C^gE7X2@_25O_]\2\<:QdC[Bb)A^GT]eaUIF/+aWAWf@O3Mf,g5OH@^]?IM
KC@?MG,6O_fCfIZZ9R5._R9_8Z+BGB-\Z(EM)#gG2.^NVe7D;PN_f++:JDI<(eZ+
XJgZ5F02#YS?_\_aT@g>0D[04/Q_8M6TZ[.CI(6cc>@X-1GZ.Z?R>82<T/LeaO_a
A>OXJ7&\g1,V#T^2K;J>]c]05YPM:d_dO?ce[:cWLM#/([USLKPDfHc6,A=eWG(K
#T2G4VS-V9XS&U8+?,GcZ+M.Of_NVJRVb;R2E(#[>^G57AC,L\8Y;b]e\DB[DC8G
S-LLN(:Cc_edKG#?+<W;a1<SFaXF&0aEeXfW5:2AL2>H<AL^E^]Kf<M)+c?#,#BP
>2:-R;NVW9[1DffDa#7?+-[5Ja93E5_S-f.]-H^=>KfNXI+AZJ<^2\=0=X8eeZ/e
46?+#0-&TNT(]3L3=8CT8c&6R,L.A2NXGeKgSKJ.Vd.SPf2BbYX7VQ0M4UIf4P1]
UE0P3<2:T/_YN?9D>&4Hd6JGP8W6HSbP@8aeA?e-]W=HM;)P[aB@J]@3UD:-4CQ#
Qa#P8;F#b^cRLa.09YA+G]99A>Y4KXV/FN\C=/Vc@M__+I[UE7)3YV9cJKYOU]+/
9N7e\U(SO5GI(CS)&DU]:]0>cfD((+^FBS\=8](:#_Q3XGK2S=IJ2cGeWV1QSGe=
b107B?=SFaP9WQa/JS,eRJg81g-A:#U5,=01Jd)U\<2.XMBg0O@a@IFNGN=-O_,S
->>5(XDRSb<c\[DITQ2g4Q5gYE,.=)FZ(V.-]V<4186;]ZI>=(gYTaeS]4G,-dC;
Q]WJV29^fE^_e.aS]Y4&f+gIaWBR]KeVX(MeI#LA2c@K&RX\&M6BS8[#gJc1U9(d
WP,I[<8H#aJ(NY+]IG4E5ZU.8F.1g\eMBE@FQ5O.T]G@d>,D[Y7IUfb60RORcEL4
_UQ^H6AK<,eUENaYHQ)d[f/d^FLfB/JSR=5caZ=J=_>/V[S52:dWMZL#K8I7-b;5
Y=-3V\bg8[]&fg9g,8X]?:(3U@=M4J/=\+R_OU.Yg>J&S)VJ5O#;,PD[][L,L/<1
1g#e^7UZ,[D0X^6g;9Ne2eSH;-cGXB7c5>AS0/5D&[)P+M8D#D;&<A_[/d4_)B[b
>-^9/[CKeN0)S7>5=PBY:ab@>8[:_SVJBJDaa^C]=5,F4@P5C^D=0^&VJ+\Je.;&
_\>d:WR(JeR=BNNObV^+6WP\+[>eQ3FIY@4:F][6g?=S8VX#(f0(b?@g^bOSa_JI
X9@TEBC&&SC,cB;Xc7S@_635(4F,b070Y>QKK=AHD[JZ^?V,B4cb&1(5a4D23I6b
O(]3OLK3E0]GV3Y+H5@2_(\O9_^;)<4;^S[YV9b)\c#,0,Z1_F2^@2@_7ED7V^@.
G])^eME)-Y&.-K^U8/<d_.-9(gB7M3N6/W\aUU#X:IJO?6?,ALU\DJ;:-7\6EMY0
IOda17TS0eJeA8(RZ-G)@ZN\fAU..IDgGP7)?)G9X7\@c:FEH.#6C0_PSRM]&<.F
N&WRF[GGD-OCPLL/<cG5b>8,2.OaO^GC<HX:_;>Y>6A41<>]5D_dLF98]K.-aRaQ
bf;=ZNdafT@)gO79U((3-H4Ie\GJ)N4;QV4Z;FfH1)KS&/QH9VdCD6QARF6d]Lee
XaeXT(d(5WX/+U]R-7T))847AB6JXMV>4]Pa<5U3T;,R6RXLHf;1J1T+=W7ZB+UP
>/^[JRSRRDeC&6ZG:;d(JROcK0RH06O9-30O+@1\aXE+5KcKe^<K+B>HTU9?G;2#
T#G,.2+Z7b>R@SH1P[[C[X+UGO#8]H,Bf]R:3GdfRS?U;RT9GeZQf_^2RAXISKb;
bd5UPCQfPB?UO&YN6CY4RDNG9^_:V&X;V-G.5D91EV5Q=LTNOOBWKLfFGO[)IC7Z
6W_L,3c]4-_MFOX?/:eQIF9g&:+If#ff-GO6J_MA7U>_K(,JON[F&5.-Gd[EHd.L
U0Q5=9fF(.KA?KP1cD689ZIQ>G&W:_F-[P.95.-e]R//HCQe8B@QS\,Y7:_Of)<=
QRI0<&./)\)O@MF=H8S9^+RRPcg[J+/4g?<_&7#OM--Ha]VV9SOE#H?4H/7(.KId
(Nc9,FDGc:d[FOUd56B:WJ/fIU(?G>U5HSJ\,b[U#8PZ42SN82_J5Ge3KA3/J@4E
VIVB#BfJ[)\YJ7O0)b8(@Y;X.X(7+@gWFJ.2LO(1JbUBCRfCS3CI7,F^+2Wfb9d]
,3g5>d+EQ<FF-/&=NZ4V[SD[e@eP+B2H+FAFed;-MPT7V3WK)C]aXFA[0SLWL5](
5,H;;S5IVd=AB:Z_?-fG<X7Ib<;8TRCS+:V4N2S.YB,&<g=SZR_43W&GZ8g_>=Da
_bVQL<)T9f+Oe1<L:M?S-KA[&H^#+^6N:CW#AgV8MMe#.L@/+OG[^6;L]@MfI#8[
GcADSADd;7:E-KIA-OKJd&VLc3;0UZ,IPf61[JO36AQWR=5>P(+S/5EN&;:U10-1
,a#g[(C7b#<SE7/g(-@2fGUb3OYe]M[1V)7/.:::<[MSL/Y76g]ccD].23J[H>3W
,-G^=:EOR-RNTA,^]a?7E/]@(Zfb0YCTVF[UP:OcO]/I-+FX_-F8>7<R4I8.;e49
_[2f9F?).N;C==<GcRA==7.5CBMcI194B.XIXR(2B6]4<(/K^+8:A9(_=LN-E5&1
HP6>@[\<>+^Ig&RbU;<:L0gW_dV12LG0:4,B7LG//a^X^A0W)L,LONGde1>,J;dJ
PPRR^CH^b\+e4-.TNfNG=+D^<4Y4R=#@b&16PNIE\#&D3Wca_)gLfBP@HUYAc-VG
W8]FF7.QY[_^<O@6J(RBD/:HE,C3c728a0&L>7/,MFL5]S)(T#&Q9:)d<6)B.B]/
VH.XOEO@a-cRF:E+E0CCfUOIL[>&DZIMTSCJ.>[7G66R=@&PF4&B]>X&L#9GD#UM
WS8IbcfC487D)QG&2[;X&a[3+.(bWHPQ(>d6P#>7LcOC9Wd[0SdZeFW8T](&QQWA
OZ2feVTVd<Z\cDOXB=-;#KSeJXJL7[4+FY.864J,SP-19/OFA-]&D@AXH30F=(9J
JDK)T=P4_8+YgV&0Q\;IB]cg=&W_SW]TSNCa(#5V7[@fXYZ]KUg;WPO/CF(:MH\]
PeUTdKX3fJ1W1HL3NLJ3XK5Z>3OS3RW\U2YQ.H8RXD_5G98W)d;NXB:NEcbW-dTa
3W&Q0C_EWXNe:7cR4\0C[F2R]JPBf:6Y+@RQXdI@IET/(@3?d9+S_&gFA8Y1W6F3
95-W7<XZe;/YGE+((9G:+d\0WfYF5c=LP&VRfW-LDa0F#bX,FV67R0&(T4\S)GJ1
b1RZgK?JY4f@,Me;0#,/Te)QdMLG(e4>2e@FX]^2P#W]];J0P^\DOYX&HcfXZZ@F
B;_WD+;b/IIJ]Y;+6EAU00&SaWRcV^4f]^^7dQ3Z6b-C3:RH0Af]O:\^Teb>90_9
1c-ebbWJ)gR]?;cQ_2&Y)55?fGC>TUTZa_D63^&S1<MTf;?(N_V+3O;b4GIgE_0/
N]D;&.Jc43E#gc9><A;LLG2VO2)IHaC-6<_X__3+.9>egF;B)DEc[5bV8d[JCb(,
Q:013H)Z,5J^DT6X+CdRcL4BeC:e+DCBLI6JZJ?17M^TK(&V8:?[=;4\K-N:914Q
69AWQeEL?0]^=C+ag_ePb=+N^EXU))F6TKC?;VOc[O-T&P8_BWXV.Aa0YbS39X@V
0>a@:TVKWA^>E;/?D.Y1THU?bXTf[#\]_;:,EX.T;?(72BO2@B:eCfH++g.g^1e8
cLW[eZ,gO)A@1.OB=9RQ3A;Wa79WSO,T4/ZY4)fd9EABHa^.#/]Uc.,I(TT,]D/9
9X+a;JZ\FK6@cU;SA8/B92,FZLA6I=RD<GR02bDY?;/-293eHAJcbC0aA(FUP&De
gQ(g4+T4P4BP0W^GXJ4V9f@0&5[6;+c5X\=8\?JAH6.d?J6g=EE-;b&ETIBeWBNP
Q?b0ZZOUW>La;>cg;>B)X8J?.Z\P=U)d]3R,@9Z5,Q:Jg_V46IFQYPFTFcbX/U<Q
#gOC7#-KXSNARg<LEPbX8/M?<XKF7;Zd6GF\c=+dL0BaLbf-eNcBI-(58+YD+eg\
K#B41X3C[FEP;[8?VeSV2d/.D0.&gWHb&F:=c2Sc=OggH5Y1]+HA9M#RFM+KKbXD
[).:6TMaX+I)>C[PI7([Kc#H:=XFNF_HEOBN0-.ZY#g[V@YdD^:FI#1XI8?J0f4H
J\eR?<4;1?+-EH2T_UQ-gTYMc^;U]S4L(?7K-N?VTS=)f_+/HaRNB3=a4BO3-_9O
DZ<EaBFScDD=P,IQEA,ZEEO+C)^8&9]R+1dK,/M/_^7<H-NYT,],>E90E_e4eK/d
7HUb_(W<;6&:D(1;fc\@;SK+GaTA25=L8JY&U)+VOXKZ[G)6PX:O-?0.>^VPUa4f
Q<=X(DPLHZK1e])<Wb#)W,.)/1eQTEJHK=dbG?^ga^58S-8gXb4&g[2U.U7#8e.0
Lc0S,R11EB+GB[^X,ffLG?LRM1Y&PBJM,_46feTF\?YbKA7@d^TPZLa\Y/XfBP&@
FYge-R2-eJK9L_X,O^I7I-OgR6V](CZ/QH76_H,E/);We/^CN+Qd_2QV1XMK[K69
TdY;2?[7cN/A5-N^>)+eBN(Y9W8.c>LDU.8ADUKC[,M;FD=V<T^[1]&12X:d-CA4
aJYRedL<LRVgH](:cDc+Cdc&-/Zf(d7>QN\Ff-f2GW,gD_dS=Ug>AQR/NTA\fZMa
KZB2fQD=9K466K1ZT^c]7QZA;cFC?NXbJ?)F2<,Re]/LFD&d,\<9:@,gdZObM).7
./]Z=,KP6YA<\a3M.RWaQ#2?Y8B=_AMI@//GUSf#g^\=_[I>)CFN:gWU0JN8L0ef
>GRR/a:2J]_:8TLaZEN3].>\;]J-\f5UORA\PNMA[8A&af5bG8F8><]EQ^1.0=PV
94-J<YZ23)7OY]#:G^UL3b;;,1O)H[#@dfZ/9>ZB_<J)e7g=YN)(#8F6,WU<5N/c
>0@9QgG.Q]2&@N&#X:6a<(H@6/0J/3.aNS=Q.c]/;;PF\>[#3/:A)fa78<aJR0UX
e1<6N7P)FagB4?FIW+_>UcaE@Y:^3A29J><)_GagAG-)<36aIFe=(f1PeQA0&OXJ
GT^652VEQAX#)+g/8S8_PR4O1HV7=Of:0)8N=>5;3(]ZK.B,/WQ,-0]#_2KVB&SL
-F^><]6CdALEeA./L,CY3^O,,F+M+5+3U)CE6@09GXEK+V[<88fBXMdUXRO]F2\L
KYd:UI=NVD9#[4TT>XAB,--(-fW^=#[?+O1Z6@fJ3J1MXc;5_J6EK0&Db#ebG[0K
Y9(^dPU:e4PXXUe6MUS<A.-CJJO6gcLH=^BHE6?4VBA>@GbZT0-VI^9^_8H^.?MQ
_R12.S<?Gd6F[;D0&1T(F-AJ.N0_,?<](<,;b7I>LA#g:.JG9P&T/1JMSc6B.<_H
Y08S/QJ3<dU/M+E&/(]d<:J7#X(e-0Tg\ZP[X]3,[8b.d#>KZDMDP-ad./8X[GVG
_)2IZ]87H\T;^(>[VUXWDd/R7WBF-b.NN8EA[/9]JeZW?:-[[GR).S[LgP[O5#U1
C=S)=-MR?1\N8)6_34Xg6ONA-/=Z3Pe7?5WM_<cTSPP5aG0U;L>Rf_SUL2CWRTHa
3S(cJ0K@e6\J#:=4f6&^(_)(/)L2UcX)Xe&N5M(I-S_\[ZKPCcEW/S:NbgJ45[cT
aGd3F45g76Sd+eLEQGW.3<eMYC(aNaAbcZ96,MK#R71+W-MA_&d;[FbFYGFE(]EG
)IL4#bfQ3I12W4/aOLN1_#cd3)O^B4K:gXB=7:U?N4bIG<</YJ+S4.[WAK9La&.U
2CIS]Q9WY\VZgcg],,b7gBbL60&876gJ,FB2QXIZfTA(X7KFP=8V[ZM@-HOSL8e_
R_J45UY>>BS]K(D:4CQ,_f2(G3G9-^..9+1,G=+;D]Z>[758F#SY7+=g&K#c\(C,
XB>)DZ1MAU,]TZ76-B0gII3V-<XCWXOS-U,JRN&Ja-UI+X?X5ECL+=B)YJ50JBDW
e704.Wg5T,V7Y<g^1KYg7XRCHKP:Y?6Z[bF\Wg7NPIQY779c7TEd:/K5X?\W=X5E
5BZ(S0ZR,^dRPCS-7(^0+Y],9ZNG>Y]/,+K]52++YS[Od(YVWc<TfZ/NP/K(=J+M
D(:6]83K;79T^N,;KLMA.0Oc1DTd\3U-AGI\CWbG)+<(AXPCTLS5afXe?Hd3aFOA
FO+^c1UAWUM^/4a&3NH_1c_aW7XUFC,aaJ(@fF^092O;)@.Q58RU3,S(T3<)XeVC
[aR@>,TE]Nb#HPV<M7.Hb;QP=A:1?MOG+TA5>4<0A0HC-9FDg1;MZ(A2\0(HQ1aW
A;D^&b_+,cfM&7;McJ.YSdC>WR_?XOe9_b52;22OV;1fI3DKV1,7^MU>9+ReTd]\
XNPX_f5<D<HaCGE[(6G,)7DLJQ\9C3Y\3Xa?GXaU/-J:eYJ\g#,>>QSNb02O2S?U
EA@UX;1[7?IX7N15ef4>_ff_E_,GF/0^O4UFO=a[1KC7Q@R2Eg#WDW,HTM#1KEKB
eR8U;.^-8K>J4[A(1?gR).fM7>@PdT,RLE:g\\W>I[,Mg;P>0JBZ\#M0RY7+HfNX
QK;B>7I:bBAc>/NggdKg2/]a=TFM)N>dT-<X_;.[>##fT3INK3W9g/#@3NNRbS&&
KdDNX<F@E^)H(F7#R38Y)c4.A+FY7.+JcSZ@HU#a2CaFCV5c@#MG=IS7Hb&IPg(g
e0>PGHHDebOId^\]0g)J6_HS9O6G/H#A&T.7NQaGdPD24:J2Y3(^LCW]F6N3I4I<
,M?dR@U#]LILcRGX4a6\&_6VI8:;?A?4KWV0.B8SH.,@^@\>/MUfH)a=1AHG]<gD
b^A6WT=^4aJD)OOe7Tb>]CZAG.e1cD?-G6#:<HZNfLWPK0+;<B954NR8S4MQU(aa
?g/Y4#X+R-(F;0E7XPWIR2I^-6C3d9?>-]=B/O#2g6>C^8L;4:bUUET?\Ra;.L+<
S,DMQ[HbHFG7_g69O@C\W:@A=:+C+Y8aD/#^TR0LOQfK#ND(A3M(P+\943dZZEVQ
R\6WTBPL3e^C1,f:=RUUK]7Gbd7c&,K=T255?/->);5cTT;WbNYJL3S1?DVL)Z,2
+;_#9F@BCKRK90B..Y3/>DWa+UZQXA=J?Y&,^G1fc:P_#>6<_AVbgR+2(62TVa>H
G=cR:E6?<0@dWE_)T=-GG4fMb;^X_8CH-[C2KW@bT[(-5,Rd=C1c;KP)N4d2C2[?
MEC)-e#SQd\3)J?\9IM&@_b7&WD?055HK)f+Yc7ZN^I@Sf3@;DY>WfX<SO,_,Y&O
[_VL&;@@?/OZ-FCb6T4<:Z(.eY5ME>ELU[f;1>9Q\eM[44F3[O#PI)8(4R/;5&^M
W^R/#@D@0>[=6S@D)7\9H9+:Eg.+^9F@\N6G/6_P7;UE]Mg_#W,3DfL(Q778OaQ,
gA[,+2L.K_SMb-]KSNRH,H;Q^G(>1<>V7PO<6L7U&V)>=2eZ]Z7\^Vf[DI)]UE^g
K3]?/=2<Tb4M;_;?)&1E39\aBP4>a70,[<?_YSg-0M;/??RW<VB@C[\O;@L_U?6_
M/fTOT=3_?Rd,627^#ST.G3cO.d?D9UHAEOY;0d\Pa2a.C[C_I5B1OVCV/QYeMTG
J;[6f7ISVZ)H/UQOAG218ebO7Se^0@XIH]P;:T8MbZe/Q7>W#a1ea^DLg=K/Y&>L
AA5ZRH(]4AOL8PaAcg&?K2Lg&0_[U[Q_dQVaZN-JL@M#&LOS2cLS8\a8,2OgeN.)
[QGHWZU<P<8NF\7Q:Ra6caNU\=X+T1^&Sf>S8)]HeGA[)cBX\3HF.R(031VSV;Z8
CK]QKSM)7\:U-;8Y]^TeMTRXM0IPL)/b0[=Q/Fc^ed6b#F;BOW78W9Q\N<9NSW)@
AH#JK;W)TN?E+L6cc;3&e)<f4O[KK.e:GO-@dR0[9OcHc.c?9L:-UA&dD].,]=IA
.V:2#8g.8Bc.J_Q2g+<,_^O92...Je4#C8dRF@6<-9@8B(U/0DY#+UF.4@^9T83a
[4b+DQ<<9\/PNY6[J@0dS_c:_JD:&9I+@U1WVR=N]6AWJ##g;9^S]XZFdXg;&.@S
0.2?V7@)f2&gIZgdC<-/7TZ_E-AAPRO&>1#C+0J7<SW8T707LUc?bO@JHEZF>Z]0
(F5SDSWRS,CR8;:8d@S56C.B7P1g(gW:S&e[3AY,PVU,O\V^g&\6/N1ccXNc6^=+
U(.]af)4P9a5IO4JPR3FE)5dfSMHLa7&@672=W2IH8FQUc]7c5+VTCN([g[REU)T
RSQP5K1d/J+SWLcdc/JOP/H=CTC:)Ef:.X>NM<C#G9bCDWK=A6;HA2&\IH+7?.-B
;QXYGg8RO+J_+BLLdfQMdRcI-N4)gL@TB:;#gEc4_MbQUFVR8RJM)=4KA?1Q7/QI
O2eMd@321^3V3M#T\_++(24Y=9>^0N^WGPaW4\Dg&Gg53GN7#_aG=9W=\;=/K)[]
f=Sed5HdO,4e0/K,.G<>R^-3;gH32A:?^X9GAL33/RPR&0]_CP5U>0dN:WV9<5P)
H>5:9E_3+I?a70GbQ+C(6#_gR3?3]eNgK_g5.8@N:YUF^84LP\J:0Q+39NPEe5]a
C0b>9DHQ4V]QA-bU1P9dJ:48ABc:OffZP@L<aAg[U.Rb[e5_R?c(gfGE>EL_QG0]
V[TE;:F6E:?f3&+169WCQ<Xc4S=Fbf2?^R,)N0WJ7DWf<A-EE<:S:Y#?c=7PeV]\
K0/@R017bSg6)LMec76HBYT#M#bO+&,bR^<./_R^/H<<8GB;&@Kd]HP4G7@H_/.,
bF4M)7KK-^P1Y,3Ld2_gZT3Ua@6^L,eQFHI9_P9\a3)IP8J3D8TDdOCF9OdY<2)g
<1=[SaLPPHV?ZfbD=>7.Y>BZ2aX1NQd:-HCRU^J[?M:d?f1ReH\UY(H/H]\FTbW7
T)\b_74]9A<DC:.OC45b,^Q=1M8EI&UE3(dO;IB6?GUBMO90IY@VPP8R63V@X1Q]
ABf)R;cU56,@T?=D@9;I9^XJ6IQK/W89dRC/@?#MbW[NUP]UA=G<3eCU.c[4SHBO
<=ACA0[+1&0=2+&=8U(B46?5f-JV(/gRa8K7[DZB8VJ9>EaI,/KG1EGdMgcT72E8
O86K\PeGHHM@5@9_d.(K&\CL1IGWfIC6ZH5_QH_5.6.6YZGbWC34L9PYW?#<Ce74
//0JQ_J0#)/5c6YVLa;3feW:V2_7P>/C/E[A(?M.WTJN:)L_5DI10F[5@@S7fALX
dN:\(/O9I_D.^dL2@Xg=0,U9,V./HOUW\KB;5De^PR>I.#OK2;fO1WaHMTZa+M&f
_E@39Vf\e7?3=O=1;(0S9-MK;;>H)QCaY#WT8]\b+DY@+e/J[W>^Bf,NC#-1#5>6
b#4b?;AGF=4_9a3<VY/6[&N[X?cB#L<?7XT_8UVcgB(D57W/?HR2-T_FLU>S)^94
^HMH0CO_[2Ade2@^_,6Hgc]F6[Y#K]N7XB5Y)^-A0W7@/2(H]4K-6fDKDTPNZIb^
4g<Z<C#&YggG]X/CMQ1Hc[Z;EKcZOSg^N0Vc4.LQB)9cQBZI2B.30WF6eR<A7I)A
Xe6Y8;9GOC?8)5=G1X@F.;SeRSV&2\5MfB3?a+AfCP=(2B6=bJP<WgZRTW@fIb=[
DXJ7XJ(Af8?G<2OT87+.@)&0H)4,fN\,NM)&\@,TGG1^Tf#Y18KMSIS[5\TGPVca
<Y\)F;5[#<M-U2^eG)_a]I/1)BG/cL0I@LD\&F)5YR_:R[0MDYb>;TK_A))YdO]H
)baE-,2(6#1@:5?@[2:;;AXUWINMaSH.-V8\FK6cI.^gQN#4d+42T\W(?T[<Hg+0
X_)4VM]E[O.9S?.=/G[PSUQX:&1CWK+N=0HUI6^g>9eZ5UMCbXW6(F?O.Tb?#6?Q
agYCGSXNA=\]cfc21HFV3+3&5IXa3eVU/AfK2.bK(Q&R+A?PPgRKLYQV.,;Zc3KC
PM[,#=J7(?e?.HB<>dMKX6=]Fg4N]V0NUM#CQSeZ?ga-1aQQ^gcR>6&fdO]0P<VV
Q4fdgcWcd?PaN(IO&=YPR)654T0?b</=dMO8S\,AH-5EW>#Z]);:1U2<8#U7MMAR
M7/]Y15TdM_-NHG;=EC+GG.c4gMW><XRZ+\X.]\>4+a>O]7;-@a,F#V:Wg_efFDI
2/(2]fW.f+gM:D^&[.W17g>a5b5a[7ZC-CWVKV>PGIKA2:]K62NM8=Z)Pf[R79\V
G-X(6,6-OH&YJOCe]N@a;,UJE\)B,<:9D[\CUZG=FH;8XVS[Ee(&&FXWAGWN;f7,
>g@^3YdY+#9]+(Fd-P_F7ZR:#5O;a55P:J(?F1=[#8<a,Z&]fTZ-:OPSU<]HY?PT
)/cWV&4?R&EcWIa<=XB:GNP&==aJc7ZQZ@]gXD@M>>^39SKK]\7cB#VaG_1.O(NM
46c/5g<Sef(<3IHJ1[9ID=5TN1C6]/ERSf2@e^Zf^]f5(R=dd<,,?2g][d0W;7\4
<APD9CCD;RAKO9b/)@H)YNa=@L+8+S?bO6R,e\&D(,V,a1IE5+,5.>A.6G[dd?^\
K^/<7;N/W=+Da63BgCN^dL7a:Y&S(59/@I8LQcES?1Y,e20gS)gA0@cQ-1f5IYBO
FIHP:\b4^<-c^(aP?YT[^KP1FT+S9(6(E<WOCE^E5H4X=8X/If_3/;,\A,--UTTe
d9GS\I2JMZKGd=I<37-de=NM48DY]U+e9OYY<0G11a)CEcMSV^5Q-d&&L)XTDW)F
70()Dg]@A2,-C;XPeNE9[1<8OM(E?:?H.K47-XH&(@C,_aR:5L7@<<_XLKaDY@OQ
JOXDTfcb;29RXP>c&7YCT18CSZH-2M4+K9_=)+YU=^6)_/M7_,)[92(B<6P.aGC8
9e:NZ3&8Q1?TAQ<TH54)99g?E?(aFcDM41@aa\g5ISd,9K;\b#]=DP,EF>=f_)PZ
T@-D(F,@)SW\.8A:[#J73[L4)D<HYGXX=URZD#L3X;B;KZ5cUGZVRS(D<.;7&B^c
W2e2U,@KeV<FQT+<\dA@S5J-?,#QPV6+BV9##P-9J<-e9WL;.2\7>,)U1&2R\5AO
7B5b=0YCUM/]7dQGd]fT(-([I-N/&5PM+SZWO[<,&/A&=^#>2,#331gM70FEYe&;
IIED^XAB91V@3JY8Of5&9Xd4ADY-W+CPUX=Z]VO@<^Q_gX#EUY3>Tf<,?+MB/e=L
F08L8U)E,d3PIB.#:f]8=TTHfRa2>UQF&A4SLHUe=Z\FSRD0[DE.8[#<.6UG[_+]
AUVG7WVYX<S:gIdR-ZI<b9PG&F)Td:9K94B(I1@4(gVRS<[9#G6OEa+,7\dHG1;S
ZT5Q+<IBUUI\I<3UI[@aO>QV6#X@+2gS#:)CfXT=8QW?f)M+OEaX:&S9C?,g>@NG
efQe:674STg5aUR+BaUYJB4H0&AN+=6D:AC/^F3[=P7IJJAYd7_^-_QU/>2(DQY&
7;@)[C[25B^:Og:@BDGbGDU8?89Ieb-F.?GJIeJX7&aQF2HM0((&-PO&4TCM?7Sg
Wb]1-HAWU#Fg8Za8bPOX<IP69DT4Lb\R1LVQV,F)<#0UY&I1dDGd1I](W=08RM]X
dF+Y<=F9X=J\ETC4;)c<AR=TA@+I.=#DMPC\aIX&Fa/U=0VQGM5RU?6??))_\6IW
YRPML-B@aa#,V3Y6/L(ZL_Z&Q7bF6HN_#?;<c1:X0d6(BZdYSIYR]:G=a@DT1g#>
S&cYHC=;R+/Ve)2AgI=.I4(2ZTY&6eQGE</AY45T-VQ49c[^H1T]d(]EB1;EW9:Z
a@HffJa\gXD)Y,ffPWBI\9B?4@3.1D21M[ZQEP[+3;^HU<-.C-TCWf9GR<81?(E=
#^N2-C;7Y6Q[@@29[^3B0:NC9c<IHA4/bPS3f=X+f#bdZ(?JK(bN(cD09^0d:8@8
X/G59;(L@0U?@>TZJJG+QWd)(;T#5d^4A+0I?-Td=5LSb57J<Pe27GYP=).75aJ(
M@DBe9-XH6RMA;f3:/4B(E_?30?(+(c6SAI1Y6edVFf0.Ze#g1GEY68Y#+WM#)0#
a68Qc_(9e6F)0X#Tf<K3Z5&WGL]S);]2^73-_LGQD/UC]:P@19+].7F[Z(D:5]9=
E7\BV?/[8^=U>7Og<6W(7GF<2-0g0N-IVc9.80b+6_TOSM9:4T6D@6G]DLIGb)=d
PcGPU[2.U.O3R^GC0UbVL#B(2gG#6\C#+CBeQY&PQV36bAX8>+6N_BL/,W6)YV_.
:ccZf:ca4T+<V_9VSV/?PUc^Y>V90a:2RLdeK;2135MBF^5Yg/@_29BCQg>2<EAY
U-;A8P;?NfKX4XKWK2@b8:#K<@6J5>1fLb[BH#V;T]UU#=Pc62/e3YcOZIWT#IR5
e?F7:I=QBG4DW;^F/<Y)\d+ed/6^V.NfPB#O?N@BVgJ8/4AT&;>,V==-9L]aO_N4
aQCaDGcO-4AUT+\HEQCTdF(SaVCP9L@E)(.#?eRZ\ggKeU357<Y?O#L(=LfISHU,
]LEgKGOEe])4F>1RM)M4&<H.U-5X>QY),Q#RMMa>-S)JVBe>VV;5&Uc^E;MRY2g/
EFM&Db#=fV-a\.9b^R;6++CJ@d0-H-PI)M;+XTgHF3Ce@&+[\HG<2WB8VdAN<VVU
\PefG#6aGO/2;)<C\UH@9&8bOg_X5NcMAeHS@>SDB3dI24D\;E3@^,2gcBB=I87f
bY0P;,dE2MN8e[;g9IdQfO]7;VIINIa,73d>7/Y?f#\05;O_,RV.[f>@&)PKd6(#
gB_),+SZ9Ig7,4BcOaI,Zb+:;5LW^GXe02L9X?KX2VIDeH/aKGG):<BUG=cURUg;
Nf)bG4ML/N7+c&Y,TKg81=(PYH\(0EAa_CU@(b0,c.+g)](>WRP\@+a)?EA[:U;.
S0V/g#I@fI7;TXWZRG7/&/)<c&09MNc_ebRIO=aJ6)ZWOO+M:C^J3KBQ4+N7KOF#
I.].@AWGN4bB&)O-a]e<R@]W?DaZ(c_@_FJE,>SHV/#6Qa^)ZEe;S9Z;gJZ#M7a(
P5<^04_8V:.:cFOJHIVba6cZ:S9&ZL#^,e^YB?;g4f3-7TJV:P6R>c^abQcWR4-K
[g]gFSRaaZX)M]cG^eO[ef<@SYU.F8_4NA_4f\Oe6:[<Kd+)K(WdJ#Q&5NO>.R\P
>18[^cL35S(&,)W^=HD[UVYXFeQ9KdXeg,&6W_E3)XcL51-QaZZFgBKZ0+>T:K&:
WO)M&Z^J(fAGQNC-A/@:YNA7aJaPUcB[eEP?f\(ECW:DZ-\S,PKQ/QO#Yd[N)VCF
b0a2T.T(Z4QYG-@)R&6MNN.G55J1X65H.XUbOb=8?fWJ#ECZ9X,B5a,;P+_FQf)/
(X9RRW?&4^a@_A6,S?Q+)fB-aVE&0W-.W8PG2&YfX.<-3<K4fgBd7Q(&Nc0>Q/6\
cJJD-&]?5GH(DcKIO7JfPMcEPUNgJeg3X^5\50Dc8Q9a_(DeAH/<L[a>c[:(I>6/
R5KdSV4BF_C.T568EX/.O.[IHJCDDX4f5_=&R32XK3,(LJIC>M2I;7:aU@<#B)J#
#RXAcG,1[MPB@&L1Hc5:fA0V1V^SMe8-\HQ;9)\U8Q2(_-H^7)D41(#cABQ;LMAJ
U,7]L9,>;,OF0B-]DGL4PLgcE0(,0<[>(VcFc5-Q@GGNcB8gScfKA<VL)QEbCJMJ
N+;<A62)_FTfQVXf7<IE6Q=?Y7148AaXG5&Mcg-X=AK/KLY6>(=UdI\WE8=WbM&Q
:-\LN78e]D[&+W[-N0UVLgV(UH:ZV7c8#K#XEZ.&?VW?RZA4b/Pg;T-19^AI3?-e
_\+Ye,#84J1RPV-5aQ2BDC0670-c1\LB-X-@<\[aK(W)WU.YA>^)JS8PZNW>EX[4
aLMMC\BDMG.)-G?AF<Y7c7_-D>\b8.C1Ne82V?.-H-E5f?UbD/YK&:a>:#UL3\#1
&]NP-acdE=OI</E6W?DfQ56fDTW9b1GSWgYc->bY<7XAAD:FKMW7DSN7b9)QG(1N
[;3[?;;D<L>Yd6U=aLVVSLYALaUQ0VZXg6/;A+3Pc/EE:NWYNJH\H>.WP8<Wec-S
>&WJd(2#aQ/J=e(?,==QJTg+MM54FKW=aV,]VSb?/7+ZX0b/Q=KXIL=G&U_JF=f+
UK12^23T\IgEP#TXg?Ge#4H/fTOXKQZ;K:2UFa[\X.:^_Y(bK^D.XM/&K=F;<(^4
?YU6W6\/HE@g37S>WGJL/;>:HeAN7#0MM8aE-eV]=26SK7D>D@N7HF[./\WF>YFZ
=+.4A0^_.OIH6Z]2X=M_d#gOcf:<D[(DDNd[^/G:+NY14-([,VV.:UXId9a/9V\.
,Z>^BW9Z3FX#ZgZI,LXbfcUX6DFO]QHMA6C8ADaW5c3Pg4;I&;(8<<U88d2NL&^>
;N-EfF,)<ZZZVJeX>B+W)A^G]VNF>S.HE4)>Ye[CPgR;E69a)9T\^E^K]EG6<@T>
T;BR2ZI+_,54K^=_(3ef_fd:<T^BW26Cb,_aD(d/QY/gFH#ZNf?\a1eA.EHX7D@Y
MW^cA0_PY0;+2CSVY)7_VX7RLgB_Xf((>8>CeS1V\aJE,+GWMe.G1D,4RT0X-2+H
TRI8.FP8JOUX,/;#MH0K,cP-;7fG\RTED;]IgOD=+M\PL?=Ye\5NH)Q(@#6FO^8&
I0B1=^)FO&H+^#6,3)H\D3:0-A]YcgS<PZP)3@gRBGQH_dIDJ0=CWW#g7BHg3_Z(
E:&a)+<[P,CJWPbg^a@70DS454)RM:V3J&-3Nd=C80gUG=?VL=b.f4c?5+>a#J&E
&2De?\)?(GCF\2F>I=;_0K9KP=fXRE1I#Mb7Ib0E)gdYZ:UI+^>E/F\b,-f6aa6g
M9TeGQ:bC3N2VZI^?G<DbcJ_9g;?8A>fQ_RbF=N69ceOB\KGBH1e65-,Ya\Y2;SE
G8]^e<H0;>WIb]R7P,^5.#(Z/_@3^/Y)50-3@-M/)3OM;[Bd2QA;CNd]\c\\)R_R
E7cUK1.f0(;G_O+1f2#:)9>WYIY@[PZ&V+POb#OGd,XeHf(#>O#XS>N()Q5KI8SD
3+,/T<_&bDN-[TdL+d2HNL(@eO6+XfebM6J)A.&B^#^a4EfK,Z+P\<K597<0ERSR
]@V)^0Hg/XHAPPYa#]:O2?PZ;@,OL[b.&:5B\M;Y3UFLRGQ[aR^RIe]Y<.?CR6Qe
>S,KeD8>\O6OeQ1/2RB8Q(DB6>G,QI+P;K8KLd:CYY//R-(XHRGG;_XANeDA(b#?
Bc(M6(U]7&E++\f+,_>:eWUfR,>gUIeF&WO@11g,X_>WFQFbVgd>LR0O9H=F/<aN
@4Y=\2^gU5&>([Q,d#9#WL?e<?f0Zd^4-SRM^RLY>[?PH:bFJ74?>#V^[4gN?AQH
G8U>>T#Ie593LL^E.RNK&2_0PfEPO:>/NNX#G3-^?-.-aS-015:dVCABB]^8bKZ>
E>3&#_Ue10JFeXOA0_d80.-KDDMeg\IQWX1<R5?=aBbSB)Z:b_5J<^Rcb_gW(Z3+
Pd>ZRH0g?6JA<L:15S=<@<..cU<b4Xg[bP+@MAW-[?5f8-?LV9:#;,Z:MJ2M9KP?
PMDHOJG^VVP_];e_6V1.FHS9-]6O]2f/CPCX0.=YX_YZ]@RfbG8B7I?bQ7SW_G=d
bBG(T8Y(UOLX(T0ef0H:2Gf1<&X8UG=f49L<^gH)/g/.MVR\CFLIV[;K\=/3^R3E
2F3YDd]D6,&b#a9GQO589,U@B1NCC3Hb>SSRD0J3Y_KHR+/&cYZF\b>-=ZL;<;HU
XH&eV.-&=FEY1T)g1UfH4X0=dRU1J)TB8I9O^9[,3T(2g4ZWA&(O8EPZb2=E>1NJ
X44&?aXgf6/JT>#+(JG1BHPD2:_H&]\\bWeL4^PFM_76c;QLL8PV&27]1J2E:KaT
,gccdb.PCC=E3C/#BfR?\_<UdVeF214SO3MY-IRf[<,@RB/QX).?1=GY3XLg9C<;
P^HT2UZI2;4)4SXADEHAO[#3/SIcDWIDgM)94JLbc@eH^;9KYORKfH6+=d3gKJO2
f5Z=3AHb;6&bVYRINQ:G4^S?b4<^S@3^4U]AggE/d.\+-85A-f&I_>b?5C1ES30Q
eXRL-<XXY.50\F9G6ZY<@4ID&J:bW,f1\;OeJ_Q>UQ-aRDY+,KfNMUfFb\1fUOJP
^_\;YdAZRH^9F:#7U5DMF[EN7-P7;FN,I(O-I/C&2SO5^ZAL6T]OUA_4Xdd[@-7C
[cGSf/b:)QP3gC,c(^aOaJJZ):d_@T:6Z_eFUcD1dWHW(R9>\:CN-_D91]QbSSSP
9OV3@V44:..aC)_4I8K2,^J=3bcG>bB]BMNM\B7A/),IaK,fM(.R4G0LRe])&2QK
K82/ZRV=0RKgZ&3eb+@5I&M#bXU;c].Z67;,41>RcF:>]I.cRaCIP6^g_?5PI^AT
SWBTNcC]J[f^)]8Y.YP=RMLF-C54=CGKSJ/CSB1fJVYE,\U1G>7<OS8WRd8\,D12
YH+M#a=)DAIL0K00_:aP14&S4>Y;],T9,<#__TB11QM@F7VMQc]:-)#KI#.QOE[P
+6LMM9eYf(PBP/Z>D&T.;fR-=a4bNS/fQKUcJV8]Jc8<+IgHdT?P/N-aWa;RA:>O
^M8e:e4DB/f3UMGZ5[?K25b#_R4057(+5O>+UAUWOQ<CJ?G&Qb9#c=NKcCD_]fMT
9fgG^LENLaaFc_VGHcgH]d,><P7CM76/LAf]7>41a5I&g5.<0)fgW7;EUH;T5La7
,.<DG.DHKA-gT5/TTZDQ2ed]71ZO8^&ecDJ021,UZ3cE)\eYYN>G)NfcR\fZOeY3
e.VS1De,WM@b=KICI?:7(A-d<;LP)0;XW^[/8D9=NP+,7EGL+=FS>#:fc;+G:K>0
;_PZYG?U?d\&5A3JeXf(N?MSQ(TWI-:cbO9ES8C5KHQ2T(W4SbJZO7HCZLA=PaS6
B5_TUYV/615/84>d/=>=STLbO@b#=cWRFA::b9+=25WgO<OD];FV9GFUXX[<eQe,
#)N&8J,(T(C:/S).1V.BY)ACb8-[7^)JYEG>;@GdXI^2>H85)=[K7PebIE:AD6W7
58#;SY##c&:]dP^Y,,e<N=M]=?RdKIR^g?IRY>W8.cFC3#Y-4aa2a3RK.57N)3CR
UQ,G1-<XYaWbK9[D:H.YPE,Vg,\BcST-e5U?[A2#/8aSeK?MCB&OB8b)#CQ[d:UT
A+5-f>28)4a0NR97)X=]IB@ZbcdTI164X8HBKd@A7IFVDU641-BcSN@R)V.gM_^f
0^=]-=QB6V9BQG?9IGGY4=?aWbK9,?0U6Y7?g2<eA2]PO]_<?aB=afG_>-]JA,_2
TX_(==D\^FNIFM4(YN/cWVYD[^BJK?g?VDg&b_)C\TXB3++I.D6@GB/0L(?+aY4N
@8/(7Z6I5gfLR9gHD;(P0_bGC-9WNIaQc:W^b\B.1)0V2Sc2=>IPFFBCc3W2@,6V
DR>>c_5[WCHE(2:5)8ZV7^g95+ef<6(Gf<?LBWXd+VD)GJOcBRP=@\YWG1CT,YPP
:JP4M9PL?A_YA+A22M5G>8:/6&2.G3eKB2?P[?0]#3NIa1\AE8(]Q4S2P0X?gSEB
6W=Z+QL&;F37YeK]]@G,-M_8X7?1<2WHdT26P3c-E=G=T1[>[5)?Q39D5<QEUN.b
aR0<H<,Q-b(9I?N#HW>8(+OZ&\2JTG14+>#.6<(4O5GL#4b0g\P<JC;8]:6d\Fg1
DN&5,5#&M]P_ec]DJ1b\9\UI0X31;\]U)2eIgD46OZfeeQeDC]HQ9X#>2-0d&JdV
2cACBK;9L94.3d^V0&BbK\0PId8,^]PL]:fb:83c+,g?Vgc9(S7_Ib<(JX\.bXb5
HMI:E_=d#C[LO.W)[E;K?RJYC]U83##\,f)AUS0FZQ#,_\8[Qf4)g#a0D:T2#g=e
?NCJ7a2>@0L1XXb>,g@Fc=eTb;aE\VO.]-]F,Uf#Sd2-JSWc9dbY.4;?6\T/+d>6
E=[5#N8S.FDab+59XTX[aWL_:ICTUTV-dGLDP_BIgBNGXU2LICMS<G1fP62&L[G+
d#g-Z&)N^2eO7OZ0RYZ>=6/>3_,1[g5&BC#/FW:N19GedSB8&016K>_e/Mb9QW2d
Lg:5eV=&^/@B)-VGWJ[.:[]G-7c239PgLg]UG(&D63ZM(E2R\Ee1657PP[Z67#Ug
Kg512=P^\&P16D@7^QMeHTaM+.)-\N_ZRJH_Z?TP(Y@/Xg#+]<WdHL/90W0PE=90
GV;68C(J8?/G;ZgZTcfg-dZ[MHFS0Cb_MZO1M^1IO]^W@CO0<cE(5La5WSe&#NQ^
7JNHBFNG[WQ\=Zd1Y3T[X^Q)>JQ7@97f+24GW,BbS);9#9TRK;HWNd/W2#HSaUWc
:dK4SMK^71G&0d7a_XMaKU@97A41\fdQ^)e0\88cA.0JE&)-:7(YD,R_<E1Q)CS-
4Ha=?-M=:De4J0)/E9[8#]1(62]B>SW9X>WE=7ZW7Ub>:I5Zd8A[Y.2>9A[L;LP.
\,T27CZ5e>HWY/SV\db#UPO\\9;c,=GLHYKMX@DYM7)M[3<1802>IO-J==B+.SOf
DBYRAW>RM.P9/E012QZB,5VQ])RJOg:\IfQ?36I.gJY]Y8#6HJ4;3V4#Q,<YL5ON
4;[_VJLD\Y-NW-H><,2+\B3W86Y6/XTe)d,\\6,6#?U2I.;d>NV582>HKa-H@MM0
>GIdT[d>edBBC@D_#7DZ>Z8<d8QLbO2e(IS[GXL0B,FfCV92=-]L+/[->)75Z(],
-Q(Ke.DE(7]>Qce_C;BS<;5Q2FPJRBH4(L8HgVA>I)g&;Ie<dF+9OK2c>A&VbIS[
gPSYC8[6Bg8.LU_@I&^f<A6e/?UZ)FJMf+bH5\+8W<c&OB/Ddb6SNgg1fC.f?D@N
PQMd>e#145G))c?a)A@(10V>7Oa55[JQ(6-:GSZ/\OZGe..U9;,,:(f83\F36S;9
GaE69W:(:0FVZ^3V@<TH2^M89S0P0Qc;#/e0UEe[+NZA3JU59TW:Y\<RT49L8e3J
/JM,PDL6gK&g.fWfGI4[;I+SX/RZ0Hf/09RE>7R[X<P&;:UeUE#F4dRZgcS+MJ-C
=_C?<ZD)V\c+]G9>W/(;3BJ1CDMUa+AIGeE-cBUZMdNEcH&bBBfWL#Yc:?NP0=H/
R(1F048RQZd=):(FO-2HMIYRf8^PVH/_U</G>+aJP]-/7],IZAHbeI9af=8ag7L[
UICfVJB61HB49)?/d.WD7ICMXUY1/6-8X:R&b_S^0#N5&aE_TW/a:GYF7N;S>bSg
1(c<L-PB[-4T7QccOa&Ba&VD.S?HU1>dbg+B#=QT#4fG+BETKP8Hc[&WM8^g[_0A
a0M<M@/K#dUYJ-J]d+[/>2H?Ga-Ya[Ff-\IeAV8JQM3RXT5Hb^,?.4BB8>MYGKXN
6XcZ8(B((fTY#1TIH_K;9gXgdYV51B\NCYQ,(169SPZX16E8-,F45K3UI#[:>I&I
2V(4FBH35#OS=H-T+68S,KLe1>82HRNLK]BX^87,aZ&Lc7>&fER\AP/^HHWTM<OI
0<M)U<bJAQ@>KYPQ[?gE_5F(X8PV5a4=359E_7NS^/GDe&]G3M3,?EdU\PM^,[TH
U3E\=+HZR:DKPd]29MKCTT63VSC.45_[O^SM1:c1&)cRa<?&^NWO.H9W->0#&X?W
.g7F2JaM/b2d/CS+X8P7R#b01KHQg(/-,J6R(CE3<VZ@0^?+1@;@T<QH_Q[f#bL\
^&,0EDI:O^EQ,CL3PT9?<,)7VHg3^\LbII3U3V^R0_TUFIf>;8ba\+f/#V^g0bIJ
E^EBJHCW(KPL)S=_9&50_e_8cVb>2_PPNee@5YLRHS2c=RZ]>,8.U\(S1OC1<[5<
9@H[NVSDQMY^fY#=1e]Q)U4&VC;MBGZDZI&Aa/5Q2E:BZ,b8#NR_H/5=M\>(HMGE
2bKIcK1#HA^BOcSO]FG^E/b1RN2XOC((_BY[M=Rc+B3UaKXb#b)X/72dKCDg=:BX
O@&503.)A[1V<37XFOHKaS^AY9e+EDbW(_dAU;_U4O)d\LXO5+#RJ+13XJD5Y=OD
5UMMPcdSM=N91G.PT?+/E5H()H-:=+?;63P?O[Qfa@J\^>39HJL)NfN&^2389](G
V]Y>^MW\@bADH69G_@S)EB(_C9QV?S^;0H4_XW-Jge&-^^16CL7>f;KU/^3YI798
dIF.5(2373DbUX83.2E&VP9,S+1T:DBe_6+5V,1@K:]YgJ]a741WP;],L<[Ie>gS
5a.aWg)UaF=CTeI&LAV-a[0YYH9)()cGE:^9J5NPWI]70X^9^P&]PbBMX0W-@]8.
J2Cb1L5O>gaFO1MCLX[3U#TEe+K,9WC_8b]#..H4aAOD6N4WD<U+4HbMdO],9;7-
V-HK]T)M^@,B?A3.KLC0?GRDe>WcD08-.14S?V9NeWB?O(KWbGSN]90[H\4#=<6A
17bN)GD+CXV^WZ>J,bQe_I9]93XT@b&8;3g/PJe(/IfVZAV;C#<W63S&RI-WCXR1
EZW@.d:a9aURM>ZFId>=4\,F(:DaO5IE9@UfLAY7/8\g>EG+2]CW@X)&KEZ/)gJd
e<U7Xb,ddTNY<(3g1XfCQ#T,N<b?E;<1@>4V.)b:f/2H+V(ZOcbKA,0g-@A5eI(f
F@.D&50J8a1A&5E_3B\0,<50eUB)OOD=E9<[IJb5ZV8T(U/I#5FL;=daNQ1Y-O?b
,?QGdbC1839Rd1eB#ZA6,E>8TfLT:A6+H/62-R>AVJ.HY9fR5J]c-O,3J10?^Ed_
S?E<16(\+RAV:JH0K;S>&1P+TaH)>Z3MRCX0d<f_/C/1DIEARe>?Bf+a-7\a\U71
KAQd_e.5KBNDcRba5:7QAGK##fY)Z1F\&;-^H/XJMOKSbAQPQ_^IYI/\I;P>EG1Y
>H&A<7YYSWab8:T5f18P)^IKA-RB5g(QH0=Jebb3F-Bf3Z8CbO97.+]MS>f6g&#7
;A3@FX,_F9a-I(:DO#0KH/1M7#bQ7./F:EHgHR([M&2]e@ZMUHRTdO#3M<,@WN^/
LZL.)3&_OHY;8XV_0cSLD]73f[d34C2H:TUO<?,)CR7cO)g,W=WARQ1SS6HI5g\J
=K_YOIDR^]RgEIIBUP<5(ZeAYb0N+bC?=@CcN(+;_98U8KBVa1W:=M0L^#c\NU-F
.4;)4#\?eLZN8+(4Gg\\c4+IBG=Fb)CMNU-c_J/T1-HSW3N1<2S8S64,YF#P9VEQ
b2E[.T+<g_T,aX1U2SJY[NVZg.e<c0ge1E6@H&()FLN=B;MeJ2S,EcSOPD>^Ue.J
2fXCe81+&g:WH]KV7<P7HB@YHZ35J,&R6cZI-8N1c>g)I..JebXe[B/F@JgYOaXR
AI;c]/fOeEYX,9+E,9P&60ZdGXBLK5SgIWMAM]Qa=Y>W[8)\L<IOaIUVVS,P+79e
,;J#4VA9:cNMDe3J1FVQ<CBWFMEe<8N]:OJM2P?1N99FXP^Pcd7+IK<,3F:_I1A^
)X&#X<9JCbP.R2JAJE&1EbYZfSf&4D)=M4L=A.2+/0(LU]KX9_NU8/.1QXZA_8/S
(2<bMV,XTH:da00S<c+_1T>E]Za2_c-7fBMa?LVAUWD/W2ITMb]3M-e;2.aLFT;.
5P95c4f27Ga([YG1(3Vb,O/Z=bZ]M(Z04PG2^D(Oc6;6Q>2IYI&(#V4OK#ZY5.gQ
X+E.H\,b?1X1-1]/&gOfX0;?@[<3&7DII?Y8R]5.[JDg^Z#C-(&b5b.Q4B5NT1WP
MP8S)3/RQBU-F_cGU;1O;\DZ;dC^P\61f<ASc_O_\@DV2-ZSJ)N0(,b-<924#=Le
_+004?5#/g/<UUESRS;8:=&])4)[#Ed_R9aT6K92;,=ddb>CDS54)\+<XN+e/N9^
IdFIf79M5K:4V@WCF#)3<RdTJBXBcWD07K5_W&3=K,2,1QJ/]&7g27<fYB&f1(/8
S]L;g?^f^TS>B+L[>GBV1;7E^+\#-,a?bCFLKQG4\UZG\E6:F7@bL76EIUF3XFVF
dQ:fZfJAG>WRCO3;]1/F:b7WD+VUcBI;g]RX;YgE=_B><MfRWT4W@R4F&21DWZKQ
:BG#_\G)?0?Z2A^XF<edg&f[SaNG]@^?[CbOgEUJcHHOQU6XY7TCWJHa3</28V98
e9N)]b+5T-]\Aa3C/^b/;Y=Qg(ZRCa3TW9d1\5BJQ7WO1P5VY=6Ng:H-_?UbX50.
N=^@@NC5LeHHfMIX_+=a:.NfdJe2gagF#f9IbR>a3;WUaE:74:+@AY185Ee[5M.F
H+g[9+aAR[[&QY70VM\SKM,^BX@E?J:XP(>Ua[21<6E:S_+C;+>K&Tb2&27\NU.d
&15X@0,M@=VD6J92C&:9M&;I/9cGPMKV:E8H1R__d6e::e>N-BW+<bHA0TJ-N\Ub
d_aU1_C+16fFZ)ELBAFaI=Ze,1TA3=1d.ZG]6((N9+2F5ISHPXE&CDAddO/D/B,2
X_]4[:e=LRLEM#G:GY,edLC/51_<A=1FDB,WK6TV>;TGJHM,+ZJH;:C^[Y\,gDT_
eN+aGc?QMB@T=X[e&aOJLgg[(6UR&,,:a)N?XMXNGg?,+/7^MLVgI&#-fI1=8+Y@
FD<_LdE(WIcH@b?@P2c65A.[eG5-NSe1#bP(E:3+(BGNc5Qc2J3YHYF\cUeX#@X?
]S/#?<PY22+^-MgD_[Q;O>UKE,K,1XMKHQ>(X_8J8PG1a+T4c;)9A7L9a],GCI&R
Hdcc)c2=cG>-TcAS;@D1_X.MMBEJTTGe+M4e2\WL6#F2NBQT?3GE;3e5@E8X-(CK
ZeL(?&?^++4B^gGIf,#(^4J_F:/8O<>e>8X+]_[<c54BT_[\dCO_7E.#ONa-)Qf1
QK2fJUR>P<+YGAg1J[;NH-.9+&-<;GR5.][6>d:UW^][3W@CbM)=F,T;/9P4/#E(
8^B1_2cCW)\J+?a]DJ<#9K^FW?fUKQ+R0G=W>_&A8>dZWH4QU68,OO#^Xa;30]JR
\3]&+_\CXJ:4\OJ6Vgb?<fafLM(b_&E#3(W;8=M(YeaTZB>.A5NTBK#cU2>aQc0?
ED@NcMH7\Z_Lb6^3>2F6Z\//H<2&c.)3P81JTIUN8Q+1Td.fQS9>&cJc<dFP<4#Z
L9g&7f4]:W?W0b\;b/+VU4X-W/?:g&FHXDH=_0S54GCBBF[).?T#cDBg;;7]W1b-
G)+M1@^?>..(44R.3@a[,a(1KB7Z?94#UG2<)&)71YKDS?VMEU4C)Na#M8__LT9P
fBM;c3#+S>g\R4DIcBJ]+SQ&EOR;dd;W2)7=,Z?U-J8VX=IP:H[@72#:979)DJB4
&QB3M5#cSP;FT:5e[[Ta8-/GZ8aZMA-a#(3YNDK(6PEZ47eNH_,eC5[VMYN^)GeN
33@^5MI5,U74(GZK62G^+/C<EQ@U7)J<cVJB4J/,H(A=8&^6V(D+=Ee?a]1:/A2U
E0+7>054,[,T?Ne45OGaM+=80ELKd\d0@Z,fQCGEegQOR;X.M^bQHV>W:0(f9XF(
2.Le>Tc^,[PJ<T&1T&RcQD2dAdE),3WD4G.4Y/.X7&W5WK7.LCB[e>:Z=,B/OFFG
I&Jb862Uf@2OSFNC.]WWgL@4O8@G/6HH1aZUVP=?d5\]F;J3E.B>f9QY3QQH+#Ce
0;86YeN&<Xf>XWVeXGKF=.HaaF_#+[<N4e&K&01G57&#(X3FP#]E\dQ1LfeW\A^7
A8:<.20FJ3@7/27J.2/4::>:VTCXI)MFS.509]/CA_DVdGY4aE&DbJE>P6-D#8YP
&4U2bTAWd;>eGa7;]1QTFYP]]d+\-:1(\.)PF^aRc?dOcHHT6)VS/2RNN)HYJYZM
O_]WB/[MC)&4VdJGDH=VOK^DScaR5X.5.S639IUCTBQ2PaMd3U+LY<B&W:&\1H,D
-DaZV5aaLJNJQSUN9>?K[fEN.1VV=D=)^D1XQGddC[3G_K6N(a7>F)a>XDKF/XV6
NQbCZSWXYQeCeBcY^-^?WXZUE2I;KD>B=Z.ZI)bLO5D.ZXHZ<9ES^e;YK;L9@Q0-
cU0&VB0?.7T8b#-;LQJcQ#e=Q5,Bg)VP\..TP^Wa]1(J>7PJRK&RYd?@96/.CWS>
N5<-<\\R>,ZcJN&BbURXN..5YWMOX>VST\\8CY[^VS>]2NLF1f,4^Oa+V3Af-E3U
C?8,OQ7-=Y4ST?->MU;1+P9AU&VA39abD/,+F4b/dVc.1g:+94BX\88^\fGS0FCA
]#)C9]fS19L\eD-&K)WC<UYT,[W=4c_N]Q#]ID&cJ^9ZRTP=VOVW3,F>::M@7WFT
BS/Y^_(PTaX_HHKb_c8Pb[5.OV/XL-fQc;(L472O8_Y+V5VIea^2)1DbFHYN>9\@
a@J^<.>#Q\S4DM\+KU>&YSPcY\#\7Kfe\HY,/aZf+&-M(Y.8dMH=[F8/VDN_:(-F
K;<CH2<LJB(Q-.1agK];)0/\.D_/O7[=WW_aFH<K]8;>KQb2bB]aTMP7,eYYQ(@?
7e6deBU/;c=:M4B.H)2IdgT/b#@+<U]HH>D[P(37f8c/U#MJafcUAb9W)cAA.f]g
ebX6Ca\[?>T2V?=/bO<?0/EGO4d_g]FWC(+MY91bEC68I8<05I_^\WcB&;R_TY#b
.,<(@)fA_#MBZ.0QF;.XL-?;2EJ]O<;;gA-RH_5D(0[#ZLZ+00X+E_19B9V+.F_O
BR1<&(5DN9N,-e^V+\>[)^P1M@4e,E9\dO9RLa.9GP;BWO^GTf1dY&)f@SH@)\_1
#=TU2IK^K1R_;N]9=EgAI,NcbNgG,.Hc(9aWRBM4E&_fF0]RZWG03S\THO.+dW6;
+L5AYfaLL\#QFfFE/I(6?6M-g+cKAE;1XAd03?RMU::87S=H+bRINP[W1,T49.^B
&8aTRI,.a[0<Y63#B994+W[-@f,C+/GJ57IP#g6CQT4ZZG=O6,M0cQLdaIOYCTM2
9?R_ff?HABc(2\X(eEf\QQfOJZ)=T@YSHIKQH3RK4aLg:c4_+XDC\Md+PH7.42:T
T+gO\HH\BPIV-7]JR>a;IaAOKSYVU;g1b7]NQP4BB)\F\#V(7#&[)SG:BN1;:70?
@.3PXR6)-M.2Y\b7>\2a8=B0W2I4eg7)NP/&B4]&H7_JJW@3R)AHUR\8/GdJg?_/
2B4WbTP:7cEA?0T;4YW6#cYgb?5d;Q06+<K-N3[25Kf^b/XK)4<&_5&D=O=,VZ\(
cKb1@GgORFBEPFTTeB#dQ3Of,\QI]I\D\J4QQ)ZT+gWVad2c-+EAPMa:eRS\RNPD
?U=;d4:MOdC@,/&2V64gXUZ4VMA;gObV=]gKe@Ba>d@(KG_:(^^C]^P-9,H/F>36
e@S6X7]6-Y/<Z=;;/8JBKAL5/R5#(7>HHR+[XG<?]c8\Hd]Ld]U-.K:5WMR9KC+I
bP_;WFH4:W4W3RB:7ee]DE/B[).S)>&EA1RSb_Q_A6Y04g:G:BcW28J6]Z(B\7/S
PYLC/)USFW1S)eLF;&aH?Q]SHfcQcBA(FMX9IH3..)F2COO:ZeD6&<dSO)7CgcZP
&GP^KQMgFYZOM<Ic<Ga,L5>gW?dd?cRJ73O;O([X3OE)99@<W@\.&<UI8S=cU,g1
ZOM,)GC\Y&#8HI\XBA/TT[,FS_aMfCFQM)BXHUBBc.Q4:[I-)_QO31W=#FC+5EL6
<Z><aV=]\=BdX&D2MP3N^D0(9\@K6&NF7PFXKQYE5AH7)?Q?S3^PC;(S@(=UPHNX
?WL=cYMEZA;C.HGOI/=3_QMPF,+8>H(7f.&Q,HQN7M(IXAU(&R@;YT6S1eYU+N]e
U[]d;>^\Pd2f)IFG:+b/2&WfIEe./5N:-EGIA;Y=4:WgL7#gEbaTOcTLX<D(L-db
,,Z(8LHK(;e,U(HT7&R5RH+JP+QTM=f6f9Bg^3C;H1V(L0Cg&DOLU@3AP_d69S]B
[XMDfI_.3fPUE-2Z#G_QYCZCeb?\-V+:X0>gB/WUfNX&XW\NB4OXe21e1X1\4YS.
P-2(F0UC-PE410&,8a_&=B><HKD-OFW2?/8.>^ZYF2-cQ=16)<WMR:8c)<SW#fG?
PZE)9GR7HBB+@e#W4,M6:V^e4bdf2\0#G)B??g,DV&7EU5a<;TM::.^,?_@AU@J9
LN<YRVNB+gOOcL9[?f-c8F00;)dU1=;UNYZbf3.]E+Ka@:QLGL/81-eCNd\-a+7C
JdJ#6[F)A2A:?d:R?G]Z/UWNg0[<Q5/B:)#P&e_[2Bcf2-O6c#8?g>>H;7>J=HPf
,T+.K]e@N2.(?8.J0CGGUFG.G.H+1=PH\/K;eTG@GE#A#4a=>X]:I-I?Z9[G=;0V
@-WQ(/f]L^3^A^#S]7]BZW?SV.TUM#R7&X>?4)[Y4.[@TIMb:/;Wb&^gPOD<-_G+
Ve;V2BYgI)M_Ag-L81JT@?Xe6;C+4_MNdVIA2=4?8eb6+.#X-4U590;EPdJ^VM.J
#M2[1<FYO>/KKQNK>-TNC3,eD#=W96a+]>MC<aU>We<E]F9.@E#P)?;TdO)7GM49
=@?_\I2_XWG?W>,cUGYV&43RS:&cAHX=V46S+W7PAb?eC9#MHJY/2C(+#P:0X/f-
A[BVC6O:8NSA>eadSf#9a4?SK]C;U\TA5XJ#AOR/aWI]UL=Zcc>bNe]V)U=La;f0
R./,4B_IGM]c<O1/:TZ)c=G<JY9M#KVFEdae[,ZJ8A((3,>FY,;bP;1<6G:Cf.C-
e>#bbcW]E,K>D_T3]L+f,0.JefdHMYXg7MT@ACA;64?bNKD12=gEM_KcY-_3-OV0
a332T&IOOMIc?3R(/dSX:J[1JYQ@LCZSH508<3+]F:6Y>04aT+?PQeZ4b[cH,G.0
MFM3b5N_LEM:@a_]7[\Y,X6B3<3(^O&HK1[H^KP]=R)34(=XJ/JDcd@6MIL1WGfT
QIc(b@2AS7G?N,6;2N#0FGUeK;[058b<.7IbB)Sd<Fe-Gb9QYCP35=S.+J#SWJJ?
\Rg6D/<V>A14CG)]A=1=^(d3K]H_@#E>I^fcC.SQcHZ0ZA^:8a/@RFd+?#-AB3+N
?WK72NVeIWgd12E1dJC]>Nd31$
`endprotected
endmodule