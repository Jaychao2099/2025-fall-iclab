//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2025 Fall
//   Lab04 Exercise		: Convolution Neural Network 
//   Author     		: Chung-Shuo Lee (damien1234568.ee13@nycu.edu.tw)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : CNN.v
//   Module Name : CNN
//   Release version : V 1.0
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`define CYCLE_TIME      45.0
`define PATTERN_NUMBER 150

module PATTERN
`protected
a]_H#KDZgY&C:_IHI=H@&U59ZcA]^egQD3eUYNGW3_Na@@50FX<C0)QTKPf25)R?
HaEQ<(NZTF3P/RZ#D,FCg1J[^/-3F9(4W>Gc9PgO_K3^,C:)E/CR(1AXc(8IW_DO
?#XOZ:B+<R^a/5]-K.2V/V@B]dM7=C4=660^8TXV-OH9^0&318US^;?B/W1W5O:]
SPHOJ_:TeT,-R6IM6;F<CK&G;],[O=6S+eBA3^fCXe4GC=UbZa+V+2U?Pa[7JcDZ
#HR9[I1BAeN]YD22fW@3cUI.9>_<>]c_1XEG9a+5C+/8FX;Oca&V;#S,&4;I74G@
.N6LT6(&.3)RLgBOFTg9Jgf>a:e6>:RH)cg2\8+#_(V&1f[H+&feg_8OaK(5CA3-
;.8/U#/dPP&>G\^[X;HZbg:KUg1)R<f+^S&,F]-(S+<SF2&\;\=6UT,,F.BaZWYW
AQV+M6L-bd75VDdRO7BOYdHeKZgIYRFe1L>fMBD2]JM/g(47G-9Z#bJ&CA)LO_TT
Sc#.)ZG0-;KNQ?ND2OJ=;g>gHZ7F\CH6W7]4f??4;JUVM/c_;g^L^^e<2EGEFFR@
;D8S),L:<g[>7g0XWS.>(S\5Y=_5&=cDfC;[AB,17_#-dYL,I0FSaF)J=OR(BY5E
E<194STY4?TcBVd7eRY?NAaK5(9LGM7L6?D(XO,cY<K4aReO@.gQ=d-HPdeeUMZ3
74;:Q9?H>\=QQP7<H].gd_@LDAQ,OEcc]2\83QFb5YU+^LU83]HKf^McLW,+gb_?
,NCUBXL0A4a\1_?&Xaefg.EA+)fPP@S9VRW<VW+JM(aB&\EY91\4?HX+JCO2DQNH
7E>6\)T6_>:D+e,P4S=PS6EC,#\#Y+O(.F0;9@=G168OVDW-5C#Re0b(2HBVF<_3
J7GQK,e/1>IA?2F#+C>>FT:AROH=[\#g4]N0<=<#gBC-)&JLTP47U?#<8gK:9dS/
3T9D]W-A7)<(:&>TJ)CbNWFNf+RR\0.C#6^W6FGfXBDbRWa7,K1&c5U8MBGQWa3a
MN[CdY1H5-cX;\+@d9O66L8[GO->#R+#)H](M00KBI\VK^)g#)X<b&Y3I1:A+@Q&
T7a=ce.FF(&#7LcTW&]E9.:FLC@dd^<P81g1YV3#IbH2P>W4KU,6Bg<RU&Z;-BR2
fQ-)3S=I2TBBVQ]#dGD5N<Wb#S._VS;K42gRa2_D?Y@H>=0ZB.<dC0:;RME+cV8>
)Dg(MUQ^Mcae.7fVG>L7B>001ZFCRI]eH49-a..;cJG^2(?8I/GA?SU<>^Lf.@d@
-P(BHY>BB@(d,/14]1/#X.)6_/A<K(NP-Y?PZC)_IeW)ZMGPSLJQX+Wb(QA&>](H
:.\>Vb5+Y+4L,I-52R/PYVa2W6@WO#DY8:eOY#0T>EBD?ff7#8_Bf7c6b@DHdaMN
\?NWUQ0TcXRIK8_BfaD_25UZZ;L?OPQdOXS_?4HM7QA_OE[Q)c+3+DQMA0fe(feK
FRDVK9Ge&e(6,;C3OG_Mb_2/.[3VL?PV[@_]<:>VCUAV&8<WW8+1g?A92c0+2.<G
X]a)]LM_H)B-P.0K-&@\,YVV]g49<F,/^#VPU5HFLA6KF)&5C)XSOe<AE]@;:3K7
d3KZ1NBCZZMGZ.^b@]C&WC<a.W<Ha#S7-4/0@4Rb5C&/d:&B4Y3\Oa]L95J=eQ2Q
dQ)-bZ(KN]+CZgWO1EPQ+7&B10S8A)/+<;8::,?:?/+A(H1BGX1<I#KB+\[K]<bX
C>bR&_,(c4F<@,+]Lbd0\<3[4Jg-f+J2X7?V;5RSb2]cRF;IQJS>:K3](M+PL)ZR
-(EK4UJ:-cS625[<\PP&17Ua(005N-A_,d@G6-NaMU>UfCbTOUBN0eW0dOW?\<:D
b#+HTcA;<>VCN[37D.;/dRGfQCV8cLYf+^M(I\d@\:NAEMO4P7+J613W?:B[,XMT
4F1/NA3+:Wa,8ZYS4NM,J^TU#;b27/N.UZ@Ea+9]cCHNbBJ\VcAHD4f4AdUBPOV4
/4G&5\(AC7bMP#g0&gE_PMI6XBWbD[YWRVTGI-df<OVGfOJ<J0-Ya5VE@<LMNEe0
aP=(I;(0aI>5A/23I0A:S?,\Y+)DCMT,JF140^W-(M7eJ#J-W:&,eM-L^d0__3@#
8cQb/c=@3TFEAHb4S@e8acf^N2ZZH7Zf5D7,fbZ[31UTXP(C)B28&17@F?>eRU>X
cJPbe>CE\W4A77JQA+bLJK0Z]X=OYL].,g=U0R4\WFQJT@QN.^\BAc87cSBKNgN2
VCP;IPO.4T)QRCJHP-.O9F_ROT5ba@EM<2-eANKED;VZ1;51H+<,Ega@g?E7^P^>
U(N<@g>KPQEbf^<E\\\MWN46\(ed5P\-^S;_U.SN[5\gGea(,HSV9XENU&ZgTXBF
e1-:EKF#a2eGBQ;C/^Z8e17=N:8&I141P&1gOV].(<9#Q\/35?a_dE.X\+&8);4P
U+=-AbNa6CM&HP[:aWK,Q@3XaJVQ3RQ6:HB;Xa?UXB+9eVU#P?1D<_\SVS+AK3>J
.Z03#Xf@2\=IL[YZ((CZ:Za96<>]5WJ^U<N;W+WP=V:O;#_B4;?WJQSTde@\Ud4E
:(ZLWQ/4C?9.Nd_bY3T2A6AGVg]E&K4^Kc_ZK>32N./2;=Cd5437:Yb<07c/WK5R
]:?3-/TU/D+8-V&FF1Q#2EV7fE&f=9a;cd)9I:9-_Q(R^J35fe?GK\Qc^7/FXBC5
4A@R?12[Wg?&Td(Wd07FZ,(L9\=,8.a<_);dQBVY8#+Jb6DbCg(@9b/M[4a<.b1K
@g_JcVR#Sa.)Qbb;bg^3-@>-/G)f\HLac(+6M\SK<OAFe?8L2d)&P<:J#<Q2HSG1
V6.>fY8[MK8S=TD9e4-[C67.b6:S?=-DY[[LOXJ)TW_5#T<L8OV-?aOFCJX3^XK[
/CDOADG.FW3E;2O,8TDN;I4A-MOV&:WdHPW)GA/:Z9bUZ&L+HBGQ@4C\:0_XC<HI
SVCK9XTFEa?>6+Q&[5SG>N+d@;-^/==Y2LAC<6[@fb.D2-#)C.L<PSW5(74>SKGg
c7DK<VZSF[VZ5g4>+P5b3O@bA,#ISae_NFK#(c_;JFY[#E[-LV7JY]]Xg<>]#<\5
8#TA8Oa)P6E);;QTY1b@MB(A[^;LP)99=0-5a4#8c-I/g0M9;L+CTRP,&>+@[0M,
)D@N8()@KTN,)9/9Y3aCRKCC,^^R[F64:297&1(N\)\AHd1]])fZ[cRTX]Z@.+cY
=N8MeL.JW?G?08UgGNGTL8M+aRXD,(.]33_7@#E?Hb>#YSBD(9L9\F/:73.U)&L#
:500<>S#MAfI0H-X+g>HSa&Q_V8=3eOGZ7WQ\4B:U??K+Od_0N_Y(:_9@#&6F_(O
2N\-2/Z>3T4#b-f9+9#FRL1D/O]A(:(202N5/)6:W2/fA=+/4JN>+ZOa16?;J]4?
G><+\>TRGWSZ+RTOG]:W;,bNR]-ZH=AFF4:[2.C:a),^QSSMdUb@)X1/#;TY)/W[
0Z9(@5S<?88QcBZI@]f)aPCZ#[&O#e3:(d)[R:VG1&c(Faa@acV&AMgb7bA8bR)W
4OSc_?Z@b0C80P:>RLQD4b=2\&X@HHXE@^V9a:TO[]S>F(Ce+_>5Q[JJfdQL\[X1
BS#aF2T0XKf^+B)4QOJP7/KE@KCd:C5e>=Q5G(c[f0S@1R3Of3;6M1MBWEHWD@8C
TQ]OTN?O]O@7+EQGS9;I@cUf43>L]@+aSDfG#RZV..\M<(3DI1XFL9H9Tfb6RU/;
e.>/4M,8N+)9JXE:gHVU7918<P;P_]KfCdC(e@\PMPAcCBSZ-2gdV>STc,Q^.#)a
3\2W4bL-0Y9.Ne\\>[1D-=W+U=1=^c)c_MER[<VY[GfJ)^</^(MEUAT\JR>aFLCM
JMG-SBG\63daIEC>Qd?J9^]D4;AHZdX3MB2B[SgS1MdN(R\aA]E)#a\ZTHOa<LT=
-X+K>54Y2@FHB>::3-WGB&OZ,Ga;E]Yd3)F90;6R-YR+K^I\]]2(64K?YG9-?8&9
L;SSQL#.IDW6,(MGQ^:XU0.Y@S^XC4K@g.N3Q>I4=Abe5FHNP<V13XR<]fTgTJ2M
dXQD=+_\/R2e+:#cQ0?XO&&;-^1a#QIM]2<-JI&W&(@Ia-)ZNDc).N<>CGOg5?QF
G[;C09S)/WW:#Z_7#gIZZW/-\,FZ;U.N_OC04_dF1IbE.:^T@GN<J31L6WRW350F
Xf^9aK&+DC8ga,7P4AB>LZF[]C^Y\:\9,?B(EDa1K=eU;FSZ;A(Y/838,R[<<fN0
@&]+8eQFKY6A[g)Z/WZQTH-ZS[c+DW1#22McF7]U^G@;f+=#4C0FH[-Qf7DY8@:&
GN9MRB)MJR,eY](4Nb0TZ,5:?BReW5=M(7I^.1Q<)a>KeIIf6J=9/<XaK@BDa2e&
Ae1^8OBJAc6]6-<.?Ec:R(K:=_MX[?0cc<LC#C0B0FV2XB;CE#:9@[aaLQ+f1?;5
F4U)9d=YC<(YPUBHH.g;W)6S,SSf0-;c_F0e9#\5VYaG\S2?KN,?I?_a8I&#\0X<
/cOS^CVO=9YF&FV^B4@^V^ZD=&^9_#);]<L7gT1@P^_a;_D4OO?;H5\KMJKe1Z[d
aM&,(+G8RNJDFa0G[9X0@N8Me]N6;ER&YUY2P@W>dZX8cX;<XBK26,.1H9M^(DKE
J0:c/UBMb=fB/Id;1C]@0GBAGS9I,(2dB@>0Y_O2:&[]ALTR5Q:CMGO?]YK,J5af
4,O52(MAbQOGIV^(=J).3KH;J6M6AP2HKQ<&;>H\H0P1]SY7N-C94V=d=1bdD\\f
61HgV=.8N[2MMf==.3X/9D_;gWBH[:^8EA2^AO1M898TLG7)TN[D>fA3>KcXeZ<L
+07LbT6\;KFI,Y/fN.Ue5;(FT220-Gf/dYAFVSL.^KYdE^CY-f3ZVdC9N^L8.EA^
f)9AffV[5U;98^R]N47]eHgf#DA9(,DXAWW:^&+@Q>(XESIHL36?0.Z+24,KVZDX
0b<)dIBK\J:_f@b4=(bfE04Q6CF4TP#H,gLO1?dF(-]=\bg>0YHdb&)eS5&1F:PC
K\gK8g@DCFd;=)3A)Y@PX[:C2@21(^\X2R#Q/ea5^f2YcW[fEK3U==1@4bY--0IY
.&g;4E]7_eR7<CYEF@JbM<J5.4/Y4Df7504^C)GLgO=@bPN=&,+eHWV7#fc_?M;G
(><(Y6@NBI\f_Vdb4R1O@Obg)Z&9>-?#L=e[;IWPCIT8F0dX;)+:WIb07>K9#-14
_BfWeg;B4E>6,#\>_4bG?HSZ_US0,)#9N53WCb@U5ZaEV0ZgXJKWD:GHGeEE:c1b
GXD1a=<OY4,6d?.CT\V8EUg2?GeMHa8_dCWb=)Gg&3^ZbO-U<4:YOA??UBNKg7)/
PBL<G/[)YVVJ-X==&>CG?<,K8@g6_TEcKAV7>PNa:YH3BR4N<([LS?>agI#9AYcO
]4L;T4,_RH1WE+M<\/dL;g)>g(7L5\fgLHISHX5b&Q\5g:7[b=UMcPEb@]91N?@(
FD6S);M88Q7N\XR8#>WHcT<8D@8fM/fEdI/N7IF@)?08=cWN/(^-+HYD.F=gX_J-
BJb9X]T5f1^eBWNF&?Q2NH1NET8c^:64fV/A15OB6I3.^;f;G[1ZDDRGZO,a9DJT
KTP9LT.4d?-US7c<IE9>bV,SaQ,XLU^7TU6;F4@V\MT#NK_MK=\]14D_LSQO8Q;6
#3TPX>RW,<,(.UVA6D,;4e.V;#TdK&bQa,d8H6[HYZb?S=@cPRP]:4OcVa[SWGYf
fEd1XZf6:7P06@8:E0_\CP-c<[JUb5dQ_D9<7JB]M_X,E]W]Q_L+T\e(19R718M\
gB@7B3XVZDf6:1Q@e<+02>[T=LA1Xa,7B^1,f.(<^a49U9I[#)/L_6=?U6GdZQ\6
V:O^MON.]CfF=V+B6D0>;YK>\,0+8)?cA\(9]ITbH9^+=N3^//:fWC)<U=1:&+<7
\K=>EUd3cN:4I\\)_d5[:,KMYbKg9E5b8F=5bK#IS\Q+3S;:+ONRf]:Q3J]QAC55
\Rb]6JOQD8=1?];5#20Ma-BIAbNW^F6Y)FQLP3G3A#ZX>A5TK70gX?90ca5;1_8X
3S;Fe@dK,5B#>.GOMZ-3:XBTbL_35?NNe::JAc\Q]@D,bN[AB^Y3=OR,e,9\;B/U
ggdbR>3e/HW^A<0PH^P_UVVLB8>2b0a2[LbVf/>B0;#WKE;fNCf/e(e&FY.g010N
<Z&JF?S+9X,d_F1T<JB)TP(D8,gESG1]<;P)UO)aX?C/P4X;/BDeFQC),Y10gBLf
M=[g)-JLX6X4Q0UZWF6Kd;6G2XfQ]-eN-:c++U(I36Qg&e2ST].<EX[gQ#W)@;D_
,\,K-1F^-LU3d0Z:<HGeOK&HR,_(?Ob_3P_T[Na-@L,W[[#d.]Y2#/<Oa+H@AU1N
X[gW[cBaMAf-2(R;A6^7agLBNC,gUZcW@3WQ<P4Og_2CJ1[3VB)46[4eJUaXA_;L
SG[DW.\-_99FRbK^MeQKPV;d.39S.JJW.g&]Z#\1(=/bJ2+.#(PX)[:Y:UORFTVO
J\aYY_YH\g.NQ>W+@FB1/[Q,D@.ADc42Y.LR.@K[c<aU\a/N7IJ5Q#KL]V9/]E5&
\MLWW9_g9aWXH1D7cU\?OdL2-68ATb8:/5TM<Z:RHfA7Z7_NbUbG>2R=+bN576Lb
E_CLC-ZJ5-;H(eb/&90D2A,4E7+Q(#_?U]]-W(Sf(#DdF[]#?@<UEaDW&&1,+?WY
eIPAG45Z5(1R.9f2)C+#NBA0\CP8dSDgOP_\=Sc>^[.XTL--S(07.9A5^T;Y7W@V
ab(/=OR-gJTM/W9;[D,7dea(IQO^?M0ff?0C#[YU/U(B</Ia?LS?]KWK#&,_\I@=
<NLYK&IA7UWL?:;5IPR&68H,Pg0]D>Q.Q9U4:46bR+93<4M<e(9b92SR]@@RfLR(
C_CTW5S4X2>W_E#YE2[HPD5)d)4H1dU8T.3cOY<R5C/c@63NTgJD&_[IB>cEX=Q,
]+W=P-P,:gHP,A#TX_0Ta,C\E?GBdK^ZE+&A1&:E<Af[++I-Y+R.5)9XC\JS^V-:
3ZbM9/_?>]U14>K8#H;:F@XQ,[f;L5?E])1,;\,FH\BLY:LS0S;R?2GGK6gecUca
(,fdNV:T#7IWA@UEd,BBXaRDf3bDd,440-f_d^4EJR?eM=aK14AS_a<>GOHJZK:E
HTO9_5KYH22SdQJ:M+JFdaP\bI-Te]bOFD?aA&J8_0Y)Z_[1I0(>PK6Qf2MK0f3_
SH7C5TPK#?]D2Ra?4g6f:+Bf?/HLDS\Q/<9>QZJO_RBgD1<N3A11#VI&a^<]\_0.
&2aH[(\YLefEa=_,?RceK=RIEKe>NZ,a,3?6N4\L3FX_Z,^;9]CS94UcXI]1[LY+
4c.2<I],c54WEFCLe8?T(M:]@>a(,6@e<47\CWPA.#=e16D+?VS+SZ3_1.cD.>J_
WQ-1HH939Q.R;V.YKOR>][Pc,S?#B^X8.G]>RXELaeMSJCUX0+6R^Fe+AO@_g]#U
g)D+GGc:gdCXZ-98;Q=LZH\I-SNG3P7./:1+U4YT2,QXJ5YAEW7<A&9(W@FCb9<P
a;P>J9g#+c9GQ+<8OHRY#?=+cB93A),<;fH3P)IE7Q4VAXZ6CI^=1CL=&<ZJJVYC
KY>OP/U9Z.PMUdQE^.9RC#]OKH6Bb2,#\2g1[bVW4;TdHMb\^RODaG)F-+Gb4JM]
2KG#E=&YaUf#?@>OO3;S+@b<&@JQL)eFGE-[]gP/KAg<51(SgT6KCMF((:e8QDYM
V>NSPG96GV5+:QS.8<A-YZc;TGE?S66>4<B#T\=E-QG&V:J?:>/Re&g6QKR37.9@
=DLRFF^HPc/gUB:W)#<LF<EDW+0.H41N0aK&6?=YcAL83Q\Fe0YEM6Xg1/JMG+R?
ae&b2f&HH8W?=]?^b@8>(;e/()[86]M#U&Rg2BTf2@O)1(IHA,[63G->3FF]J]^[
M+R;2T897b-W?7SX>-d(6@?E1e(F8K=IScb)\V./@]_\N<DJ6<I,9MfP2:,OV>]#
?-BJ;\\D7B+O.LD+2+g8[2fUeJA/I=#P3W3W/6(I7V.AcQ+/OMZVZGIb&J_Y3_7g
)4BTYOeAV@CJPeFU;Y8f&C?\F/Z&AcN(V(I4UHMR:?QG[d57TB^@XI4RbdZ@C]43
VRUUJ/f[HT>PWP3c0#Q5Ve;]U70)E&Q^-NCCNWGZMDBFeNfSg7XH17FI=bUdc]P.
T2U<O-=Y8\deV[1^@P>)QXJ6ZAN[U3J:OCCKI_1A/JJ+UU\1f;EG^6U<OQa4JA1@
C]2+a[dYJfKfg8)OSeI#Y.N/9@.2R:,O=Gd(gT:N[6ISA?EaT.-.BPJ#HT8SXBY=
3<;DFL.a4C9:>@=Qd=6c.,H?],+PcPL/>V\<AO:]TZGc+LY#7^TEE)2O-9_eFe:G
a<<;g[2U438g=18K>J1+Z2HE-MC6ZA=Y^MU-5]#Ueac9VIb_>BI.E)^AF+U0YJKK
fW)8-=@.ZONH-OC&<A[5RINS&.@F_MX)03,1&-@UKGdW7=TTRGU1?f3ZN@R(^b]Q
@?52D<c9^FcBe-,4S/EB.eSP5ASGNH>V668<DH03@#ES6gfeL<HSODJ=?O\O4&e2
OUGHG09-P+a&gdc-52EN09+^2IPRY^3X^J(^IgZE4c411,NYR,^a<)8EI+I5=_L@
)=g8)YKHYW6Y1;P[a7W[D[CA&JACZ26^G&5cW#-(O89A8J2\e_4AUE1GMPKbE)7D
EF5XFMXG,47eH&bTVWDBKG/O.dY+<+ZN4OcYVQaUf5QKTZ@Uf)E,3Q(IGW[e;2\V
<39.N+),?-LM-+@EL8@)+^=O_Y4,:;P+?Ob;[E^>_SgI>ZdY5G>Z8A.2.PN?L8^?
SCXIWC9<\2gJ?e7@NdEY#+a-7cMOBc<Udg3-eKE]4gCWLD2?bg1-[.c83JB/OH4J
RLd,?:&VUQ3RVNBWHV7H^8LW?3]A\Z<Q.g;RG3HEQY/Z<]?_B@Bf6ZM35e#:_-+)
dA-D_VZ,-/X0X9+:[:\00_:[TL;-ZJ-e@N(](S(E^cL75C.>gQ+N5H2N8.gU)fQ^
c2E;,[cDK:E437X;L.6P3QS53)0^IdfYQD;f/<JDQ-XX##f#M.6C=<.Y87g?YG0<
AY2X\-^36W-XT_g1:B&DEf.0[&1@MP?[NLY.LTHYX_?^=A1S=OTT_(.>=S9G13c\
<V5EF9=WYDTT#Xa7_)5]C?>_[UdVVW]LZ9@QOc5H:Z_&)C6KR9[2YFWH0=G#:4Y9
Qbe&a]^>GIS7_HV(FDNFKMW?bQ]C\N(2>X_YObG7[SQFZecQ1gG7<0]8EIbG?ZGE
3Id?^eRe.LYZ_,_]((cN+M4YPe:LWDBJC;DW6#,U]Gg.Tae2ZcTa#^7Z1YP-F9MD
]SHcS0^-@@R800;#DDe2Ea]V/Id)FD>dAXZ./TeWG(:a4Kg]^9KUD11666eLC/Zf
VNW4-Lc=NS8B^_A+2]ZL;;@W+SG_KJ;L]8_1YJFB(BJ;HG^B4VS;]-cKG:b>@+<L
R^GN@K[<GQ7;U7gW^fBP<c0G@fF]+SRHg-/KT=IIb=VW@eL<FN61V+YCM#16;)XG
/2I>:K_-3P;H;VU1VGE.ALZE^0CQU9AF[^:77U>fS5eXYf1+7177@BF9N-PfT[7b
f@M5)O##97V8A1+KNT2KRND<]R806J39#2LFe^@P&>I<):1G89c-5RSeFLU#OLBJ
ZC6N5VJQ\6WUa5SHTKRBaEPU\)^@7[_3,.&VEH(8JIH8M[/._L_(>;I-#.Fc>Rff
+]Sb-)0SU5#e-+63G+P\ULd?:De6US#Z[1G#-USI..Q?-\.N\-EHW7I.IC4-M)1H
KX2OVeK8/Uf@=T9;>:-VHF/+;^?KCd./PP4+c^J,[_T25]C/&D&gZV(,<+)\7MJ9
-82&e/Q@D2/Ia0[\9(>+a=B(#S0B3UX<_e;5NedcF9Fa:bV5FBbU:M11G)H(?ZG3
\KA3+1NGGCEO=WH1[g0D[X<D7^3<X<fX3]V;PD1&E8a^[_FXTdG3@Q&>@OT5N3=O
d_\Sb6eCfb:)8JY;f>04eAP#OR/KMXK/g)W-@/QCdPRfbQGHK4G?JB)G7]<KVNPD
g+B0:WTc^GdE-AI^8W:4#]d28(VMJ=-GG7)PJ-;Ec\W(6a^W5:Z<4.3L3/=M5_LW
:2V8Q_/4PDWCbNeC[B7aAG.Z^W,F>1a(5bY<;1\4[?)4U^D6]Xgb.TF34bg#44bQ
0EOFS7^W3]RM^6/?4U5Y_VK8;LB-)\.K[Z5\VTbdf]W?dB#8QZ.V-G0;N-,-D?Te
5>//c2KSN.eQ\VIdD3=M:=:V:E1Sg9];-fI(M3-J?9^;CaD#<H\;Q186NKKAZQ,P
\aES&NLaDIK/)_N3<4)F3##]/>U\BVL3W5Hc?/T-48<H(;A7dRH2YQ_[/[#gE)?I
EE#9=C644aUCSd,9&X-,K2-VRRSIHR5e;E3^&]]f,2,^9[2e0?ZDQ>[N7&&3:Z0>
2;.bE^EcG08aIAbV0eTE;39ECOZQ26FXCTP@-b?UG)5F9M@eG9dA;3VPZKPfJAa)
?We/-_=8^T](O&6;_/])MZ&N]eF(#PQO,5gNe\]f[>&>&bE[2R+ZR1_IW/A)8C?X
2T;R:eaM>D?@G93+DDZHb82PCQ,&M<9TG69dQGb\-NOS85QT):+/)-Z_5@9P?^)[
N\KA8fB1\0-[(>8Fe&]^RgP/&CV__VIdR(KHAVU,3>DT[B],1a<Ib-)S4HS@4c29
E[7QRdZCaHb[1.X[0g@]RIHgM&+I/)&;87aU4[Wg5,XE5a>=fK#\B-37GIZOcF.9
BRe]1,ag[1=-6.84=6@@7gT]eQ63/^92<KJC0-K_(aM,5]VaY;TL=68PXWe64@#W
YEB^aB//g_@?F@aMG8dM.CDJ\W10)Y]#Q6:8TLX(;&V;3<f_MX40QI[WJM1T,[8A
1D71J?.0N>Ce,A&A8afR=)g(fb[f^Q/bECeFad3@HFC\6W1CLEG)1VE^Iaa\:[c2
[;2U;e+M-b2Z&QfD[dT[4=GVV@O,/bI[HKM+e;F>W>P<B_3-/&La#5PRaeQB4b0.
SD2S>;K/E2f1SA-Z-9W,c<b5?+\UIT;c?AI:K@/GB>5SESGdC@aIS,ESRcOd<6_7
PA.R@7gT(UGL3/^F?.+O1R>?Y5TL9;>?N@-/,,.D?\(_,\]bS]K<BYZO-R_8K?=A
M^K71Z.IRYM1/IXDPMdF0^MAfY-]?)J)NU[VP3(V)8e@D#ET^PdDPXLA4JgD0[eK
/bY)7.XHH6I(;<;1RQ[=M&9N@?,69)DW9L&1g8fcKDUY-)EgIG9a=U]&A1gH5eeI
L>2-bGb+R5FGE=;H\e;d8H.:>O1cB5B_0^SfC-GI;)OOSA(dVTb;PNXV@dL3;a@D
)=IFWf>Yg#b_/=-&b^8&9H=f?V(QYM/HbcNS4?KHSG&5&/ge[6E6=74cKUCe]cW;
RW6TOFVfY_0KS5W(4aPJWA4Ed(L/(DPU^OTDFRNdbB9UVag=g#+A2@H\aRBTMOEY
;:.P[L)df)IQ<3DUFVRC?c9c/9B)=.([Bc_L.S8N-SO7)QO1]CT&@X5ZcU(<T=Nf
Q96N;:[J;BTZ/.EE)NX;VCH>SJ)_D/HE2T[eY=HILCX&8;b.5Y;0;\_g,>bQ6Z0#
).N>Qbg/da\Jd]0\<#HegIH.MXK1,0&Q;8aP+_0>KXP.A1]I7CQM6INI;fd+Q3-O
MH;F<<)RG@8JNOKF;_=C860PX_:_B9C9]8-;UIW8UQ&SDUU,@>g\C)?8BbX8Aa\W
BEQAg>Zd:G^b2D2/?PONa+D/KA;]dZ;A\>>U:X^a1QCL1[eUUGH]Xb2H-4=C-J-[
dNAgYD>0O/[cTMY(1K&NXLL-W^^0fZI3GJ@Z4I8\_-_67UN7U9:_JO^DgDB7B=]5
>gV<TMXf7O7(^9DK0T.R1D@E1Y(HU_Q9XRf@SdU^/+DNHCO6;D7N<?HCORL?VN79
[RbVeObR42f7PH3@Wd[OFH2b-K)8NN^;@BQK[8MR&EPHWIeJ>QY,,)=UMG^6JKD=
/T7+e&;7+H7PL/5EBB9YJJ^4B544\F3+HY+8.KAQ10:0);.RDF2Bf>fdP26gWD#@
1Qb:1(#<]G6==_62L,^)RaPK24FWeI\DZ:_IX(N?KO8aP=#,V3O7O@+N]c>2V(\-
]8Z>4)(c(9CNfdWa5C>(]JPAIYOS+G&AZD6QfHA_4M9DdU[8Q\[bEPVXKO=&1C(V
gLQf/+8:#^C_7=]49=Fc<Bc>N&[a^ZQOI6_>[^\^+3EW=9^R[3gE-C#J&@BLP&)G
C<=5<+=OW89H8IBYbd.CDF@\J3L0+cIJ_JS^[BF[(Q48M<2D8=e.J1B\^<bCf@B/
57fSNKO2<gLeYd;K0/&)<bZ0O1G<Zf:N#c_=1eLXCB=F4ZTR<KEUd4[PdCF(I[I:
E1&O<SZ_0,F/D9&817M)=BH.6f9))J9)T3?P^EQGR;KT[60WUOYT@@bXIYNYJ;+[
(f(4[/d\fNQA#)WAPeYf+DTA#LAS<U&A:bSE6H.10/4:CQceg7G?O:+R?8&:P+2T
#GV2I2F(C<5[4GN=+1I](.VeXX.K-#gN\J(:QCY5X8R(_;HYL(FZN5YS/EKPH/.,
_dO.C>V((bJ)YV1&#0[<CRXeL9:b9WVVC-[.H5VMWg(#;3Q62^+W/Z?]8XO_.U(,
FDI^Ag_,&OVFXWWJ^e^D-KdW7:Z,._(_S<KGKDW7<ad\/T)XH(#;?A&GXA2V:fU-
0bfeXQ0:0D_M73/SU@<:Y]XY>1CPe^/L&MReECbEL/\PQ_e-R/Nb0FH.THfF4>C)
fUgePA:^BMeHG8&Feb-O0Z:K<8M0YbD?c]35_X@J._5BH7Va#J)EX,T9MdJ+:e7@
\)]:]ZE7Wf@g0N5XJGUVEV6D>^dL,UC4fAA(Y/70dcV8JB1]1d0:[9(P>H]5\b7K
GP^e.bU<cGSL5U#[Ze5GD^cG81A5O>9[J6B(B=T-LXHLUe)_<C_Y,_+&@R).RL]_
3S,Mg+H4_<K3I3(6Ad/25U\MNe7]Ne6U]02.(]PT34LFPWEF^X44X3dGE3aD\P,<
-85]G3:,:dOZ(Sd5B,)dV8S3M99,Z^\>2CE,((U<0/6W-QKH(Q5Pa6ce.6YW23^#
]P(=>K^f[[/[-(9@6Y.Df9Q3AQ#X::7W:CGW15](<d5]4\LII:A2X)Q0(].a1c>L
e5EMS/0-AG4<e1f]@)A&dOG79ag-RbL;GVYCC4])I&0&]#DTTaW(G=&T^A+CRbg6
]+3Bc+)2>0<Z(N^^RJ^PXgIMUT4E-F_MM84@+_L8[5O2GC9-)OdHVX[R@2O(WJcZ
CM;fWY.BH2#>@><YM4YY4;F.6QY/b)Ug.1Z+1TADOcX5>+Ycd[GL(J=SeAIIZb&/
I&:;Xg)<0JbX>b>H=6J=_:E,73#)@;e^;2-#c0gO[I0G1Q/5_K4deJG[?O4bJ5:6
I.e31JO+QDa8g)=BRL:0M/;BMTW@Y7C\YYL;f2G,YP0P5ADaE2?,dP1#V,MA>=>M
D\CFYZL?;CGG;:P,f\aUa0.Q:0;:@0[#@?>aIOcMU)HB[PcbW=gTG(D#&[H^AP9@
7P_8ENHa(.(Cg3JgUX?T.SV/g(]QA?(S3:/@FUDR@)Nfgd#7CR9XfW=7[.+GNSHX
>H=R<^1SV8#dXObZ\37UV+6>RCOLC6+fR[9FNg275A,cOYdG,N(T>E^=O#g<>M6H
^E49bd>65DSU-d/=8V.INBJ)FTRFI+>+9YgM_+;A,fJCZO\bYH\#1gR^;O;QZCM^
XU(SeDBdXPNgAXc<C-6TAH4MWW#+&HUU:ce;S#Q0+g5OR._]/#YX]0)-L4MLGNbK
--;#J:8DO&03KJ+FPIK<SHD1H[C#69DY7)72RfLDMad0]H0(S+QV9PTT;5b35?-/
984?,=)FB&51_VM0.7dV>68f\>c4<2aS]NQ/T1,.H9-VCa6MUQT8a6_41A2HLYd+
O<3OF\^.5S]GeH5S+aMKC;\E7M/Z:[]2-2GM/I37C]_2g_^ef@f-,C)/EYCLMD==
L=P53X+V@/VAJS5>+6VGac=6U#/56D1:\dQNC5eO<#\W#U&^2=bV;&11B&R&0/7\
3HACb6\)P2;X<e+F01ceX.Ib)FL,5I-3c_GP+J?T:+3?NT1=&1V2b1d>2bN9YGH/
B7MLL+,,>><YVULRD8AKf=5b)-W]<XZ9\>cKAQ&NZH#:6/V8F81RW>B]GVd?0/gY
X&,W1CZ7b<]\0K(b0f0g8BKHOK[2)N4TH[46?fWd7FT3&#\)01Oa8L1^QL9V3(GC
A5)]e(aUHT4:.a[Ref.\@GGDW64FH>QI,)#(Vg1WHMK>\MVHYL><&e#:d,a.M7\O
4F??KBMbfS_+_SB)+:17^&aXN(b=GB9_]R1SDFAQWLWg?A4W?ff/LZ(R)7H2H08,
MC2,AfE1\?<D,9J5R<Ne&XULa[+C;gBQI@WGKA.T9K-P);_AYW=D.A_,>3DNF8DO
4H.bD3.9GL0,6E^9L7ELe./:.Wc;P,NgZ6PXF---OV=&D^2K49KV?FI#SQA9_\:\
/5H?CB#-3G\EYA=FH5:J1TC^_<[b/:VJe9^@0f+CW0>Z]RLL.1SFV:JU.YV4CO.@
;]7),C0:)MHY8J3OW5dePfMS?>7[:ASTQBS6NE6[E/T&6]?RDa_Yg@7[T,I<+ddI
E6_bFNRKL?THI\#:)Jd>QOTb0BZ6M=U-0dYR<eVA5EVfWdaXe/=V7>/@ggK_aA#<
cN\7P?+EE=K)5c)cX]F/HM^UHZ<U9S;87bVB:N\EM?ATFYEVN#2L\,621JTJ@]6a
#EbG5&)NCAK7e;JdA^[]^;\#NP7P_6]1Q.7O&,L;OHXdJW_UKD]eJO_;>a+IGX>O
\&6NO@CJ80dDWcTbVCfZRc^Ma>53#HH_)49,,W6:9ED]V,a_[#+[V5?cd,O,7627
;.]gR6AJeA-AD7R\D#/CJgX:DZdL6-;cZSUgKC0C2FG0L,WM96(DY8g)?a-0Ya=O
Mec/(d>ZV8g[K^b^Ja5U+49_#-fD>,4bSDAMP/N.=E)/4+O(1XZ/RY8OJ9XU)WgI
eG[\(9MGKe;V;D3DBD_F0IY.I1+@P^(g:>M23PUbZb;KS]XV<?;)F:IMb;Fb<aIQ
26V3&Q/-RGbTXdDdRLHNbFU0,SEI=4MQcYB<K<)WB\,7Bg_;,?VWW56g0/K,.fcT
JZNX@KR_N-N(8OBWAKPG?B6&LO-?.H_@1W9AL>43&GF6;]f\-N<@F15API8JE\US
dB\Ke4bXMJFI(aD_P_IW,0eW>P[GN\-B+Ce/2[=)JD4aH>@UJIG&=;4Xg4<^ESO,
6V>#5QU1BXR-^7V\YN2X@BYDb^6/P?G<2SNUcGZN\-Obd\+#a_PU1GTC;7/I8N;\
^PKMeUW6c&9BQIUcTd+X.1/30S7K28A7^5-7J8\57RgI,e-9JeF=7F,GUIOB734.
ZAS/b:E/?ga6g/,V)S-@/0R[05SS4A\KY,JEZN]=ea-.G]OI(:_E4Lc-Y>?F&/<R
Ba9\RfUPP0#P1M#2U+f1BD4R;+4e&Kd6D,,F5+>D&^QN4[?@E@gZ9g1(B2U(Y<HP
)RSU^<1>VeXfCXB(?.GF5C&Z@&(4T.DU4@Og,GT=PLVEceXf[H?4C.TU^W#?a4G,
3C2^GWS5fQf_NK8ERR<1,4\1DY_eLeZWb26P+^>7SHK>^.(-#L@/O3Hg8ZTQK<[F
VcUDb_+XL4gc92\TRA-T]5\#15]7<,_ACK+f+]g&Q(b@OgRV;833b<]Dd>31LP^]
Z6A1P:0V)L=I0C>2fJK<-L4N]_1HVE8EV0Id^3gC0&FdJ#>>T<RF6+O2#R@0B-BL
[GdX^I3M(ZRaB(.-SF/Z9TI9@U0L9_\>4[YF1QW[QQ#V.<LL7(VbdgV0ZG8RQ.NS
/#1[@IfZ;6+P)K1Q0HOL,0M=R36P6.T:]9H227LYF)QYXd7a2<5ZKP#E/#A[dQ]D
Zb=(QZLWS;G>M1K+aXEK91^P&8eEb0(+bX.XBNZ05aV6D,47f73c#>2KVf^]33,Q
@4VL9,I8JB&>a(//A3@3C_(Te6RM.P4;A]FA8^,RP;<615,NaWcbGGD;c?B:>G?J
W4U-TMUg_>O(0<SE)7VY>[(L=MCK4Sf4V7d49a.&dQ1QVG;,+WP99O[P5)48Q\c(
412bX;,.WPgH;YXZ8eH[:N#TZ#f>J8A#T:+8N@_[/^+-?7a@A7Je<3W?3LbWOdEA
M4OReIGcFL<O7ARC9\1ES7VJ24:28_5Z.G##e-XC/5JR-R3F(Y3+I9&EbVe/D/e(
1+N@AJM?a#e9,.;^\I<KQEG]YY6UF:5+=B+SI]Q\QHMcI+5Nb7D:(JUTA>=L>_f&
4:GBWd&G&NX_aA88F:Nd;#33.^9NTN=ZaU[A;(aM68.S>aeD3/M1&9_UWR8S_?W9
OLPH8Ve?,_E#I,7f31:@/A5e6b#;;]]b6F(/QYgeLHE(J:]#@e0TN?c)\K.?O#A;
P;;E8IDCCX^B^6(e.6A<=@J.Ta:+9_[I#48>78b)4+VQQ7cI0#>B(E#.6J(;0Y6L
&cUdKO.PFVDO^0Y68&HE<G8==KC23]QG@2].2[\92T#?9LDT[]2cBQf4Q;W?FaJc
9S1_XebS:0f0W/AQBDQW]?9cbIgC0e15eMD+:<YXD@H,gHM4LK,H3_-H=K=L9NS8
ZLK4eMK@cQ[-f#EWU#MBXQ(S4.Gb=ddaJMF(@_\-:41bdT[G6]J>gFF,B05<,K>B
ZUJUH;(FMgT6C@c#3DIS^JUSOY/:]RbGfAC_d_Id.Sd?6..g2M>ddE8M?DX[6-3T
_&:812YICMZg4Y=gQf(H313;O/-#SCaZ_7;HO2V8TJ02=bM&&>A-G]<?Z^VXXA9P
+9[+8->eCNXZ<g-;:6,F+A/O;(2@C0[;39R>CQ7O.)SMA=4@]Z1&]:&QA>I=T:VJ
4/0KSG;O?(O74e6+MWJP0NF2<e1g4De>#ZKF0SIYJb\&./MC=ME3.&4I<LcW+fTK
Z0bRZS=AK0;eWT/eCNYXK,H&SG@5K,V4BI+6O>(W>\ePRQ8A7+aT;2gdU=\_9F^C
-Z_#a\5&#C.YY7D9SA[=-baL66?2Q6SB1G[+=D.cU?O9A=]8NUQAUPI[aC]aSIVA
eJ\24DX_59f,V&(V9AQ]B\-b?fdaA9eF7:N,ddd2AePVUK0a4UNH:&Y(<?;<C&+(
U;R+fE?J<AISVGZX9fJaE@:6,62SM>41=R=6,eGTF&UHbV)3Q;L?ea6L])Q7ZccI
gc(c/2S>J5W[:_3)I4fS<9?Z)Q-#GSZ2@;dC)HM\aS/>K\^Q,[KI0^bG#/G07[cT
a:gM<?&A2eVB3/],V:,MSSLB/)&2;@CQX0:R78QFgAgAB\)1Q^2)O_UDMI;+c9MQ
W?c9L0,d\gL<D51#e_;1)d^9PC0LH<_.D_M4Rc;:D@GH;M^DAZbBe)1D@0E5+-GE
H,Y3L_<[^C0BF7_Y[0,K9FOPeJIf8AYDBZ>MbBB[2^/e291X9G;].dBcM>:6Q6?L
_1FKdR3Qa#:,09_Df(EgW@F):LM:]QUY95g1\<XKH45H9GfC/H[&U1C@Z7IFca\W
HFO5=GaF[1_U&3O?cfKcJY59SCJ486D3eeLJde\#D[R;7JQ#?^@46F0#A7&NOO^b
-X6JP^bJ[3_2.aXR?eg:DbF.G^bPU.LUg&Q=/LWO2eK_>9LF^bM+;XEF,26R@9&H
,D3)]67(X+@P1f\W1a8RPYX^LH@H?7&gC0S\]-]^7&T^/X.<QF>/I+f0#_)+.?QB
2FgLDC5bEfQAJ]JSca5]\]1=(f4/7OcQfD2I=Ce?@PMQAJc-1:(_g?<0ZGQVH?G:
EMdCQ+8D^VU/ZTfW#2ZTB/QC#^G#+L,,ZU5S0+B/M3a13Q#fPX36S4bDRV(\e,B@
6QZ)b^/WW#f9U?2Ve1WU\FT656OeT<5eCEe2[Z#[Q[g>>KM)B20A01,#c-U&6ILV
OR@OGGa9R6TB1D9D\d57]THP6&+3=.AUYW]P)E)Z,<^IF^F@/c8P9A:/@WO;FT)D
]LTSW76:54:XV/4BXTU?V_^6;d&^3^@>T:)<g2Y5U]PG77)VQ\HL3]VKB,^PPJKS
.]N\&9@YVBT^XEW,@g6f2MRc0/f:2dRIgVEHV@UU4UUL:gaR4)1eH7EQC5(UM7U8
e:\K-O.4Be[.H&(#YK7Rb3];OV(3V:Sg0b)8+C^IZ/&8K76,g:Jb)Q61ATKQ-Qb[
f?F]V^]<ce@@@b>O>+XM9JI]beN/64DW2_N=W>+UP>_O-HVHQZI=^=faa<W]cbfG
[?-KPc.8NTGCMDSH,@7P_@N;afJXd9..C;MR+_QR7\R>KP499H0M-YN^SG33>Bb(
VG\MPPIaEH_368)__1Ja:Va+OK(U6:-J_TL3>:D-VR[V498W8UQb\g#eQf\N/;/S
AX0Y1)/Y3:A@:3ON)#gRd)M=68KK.7bCV/&Q,I4Q9aVI:/8eLU\ZUX<g)ODCEE[&
ce#dfSH;(Ee9)23(gP49:0YP2+&ff&6f3F9_;:1>8C;b#G)bT0/KQ^&T/#69BE@G
gO4;CHGb,D^[Hg/\3E@;eJ\V22XeP]>[G<R(e06)-6c&T>8P2H)X7eYND6I^4)Y[
dGG4L-6FMUD9@,8e:CL+&JVQeO-4MQB)I&LKg4a4<\3P4QKWZ@-2]90KN2De3VJK
/H>X(gQ/1_d3&QfD,012&g>-55AT:[ZKR7=PD-M6_=\TI=EcRFF5;6R@R83@73A-
?fb(\V:L4Y)ULd2)g#+V?)<M^@7UV#b4>O3\6V@YURJC]QIJ[_ECM.KDR2&+Y_aF
P3N+fg5Z2VJX\(OZ,6gWYHWO_D?^WDX+@ZC=R:0-J3F#@dG@I_68e+EV#A]X08PV
XKUbdIAO+4E/S6XfZS[&aPZ.2aQOR/F[2#P:_.a0[WIOE#VWAW[/>D@06/E:4@KI
;INX9DSX#dB,5@Ja5Dgd3)gJ@DC.7GP]#QASYZF:g-F\CTg5aDS6,R#ba)M\3P6c
?)>Z;g-7d&:;;AH?#84g3U@^1aA11RMADdILE;.daH>&N?Z&&@O,UAWGGbf]C],]
E@X8I].da>3[TRPb^I<@(dD&I_B4CH9RV[:BEaHH(+>[@08+4M[>Ga&>\YIK>NA5
(26EAP5g35e\9YA;7FE;Q@ES,LZ\J<..MBY8DK^ZR@1E;?=423QR:<GQL9FN&KGL
4X,;4/]/2T6BYWL_^ac>(N)/?87H.=RBaad.4L<Q1=26<N(N7MY4BI.@BKb5W63,
MUcIG16cT\bO(.[X3)20QHF:=YIBR:_I@\;5,56X(cKAXP]@8QOE9HR4G1EV/31e
D38<1<aF.RA##8Bg1,.-eM7><46MdOX\@BJ>W#eg86&a?HG<G,B7OLSeS102C=F/
.N?_8-KdgFUT9.+SWJ3[,3&e^LF4\aEO;d)M-GRVLD>@C.3G,D2VY,0>SdMJ#,c+
J7EOI41bE+6#[/))DW_+AH\2U?Q6L3Q@OQ8W+Rf+\YBB5^+2#]b732.LdD8McN:&
WC@(^>L=2D(QROUQ5W&YTcVI>8EGO5B=7HL,6Y4F;b.ceaNf#H;0Ddg[UfPg,5.)
Y;]NEBB2cSZG,F@_GJM@6[R50U7+V.cQ+C#RJP#Y9YNDO)D?YA\WG27dM=HOd]b9
O6#g(MR:I>dNC1e\Tc/0=eI6&S6JR7R+:[18E@f:3N+e0(eY<SP@]@[>WQHK^UG9
G&.XT1d&]8E_;7KU\eT[KO_)L-FPb-^.DAN[\b;@JO)\EK@+O4,HS=C[H]Z02P9=
B1EFTHKN3HE+N&?GAC)aE:UBC(ZY5ffF#6GQ92RMNI8ZB6,E=R+]a]^89#0bc\6f
FZ@+M3,SJ,0HR6g?e(H#1P^fcU;J.dOGMdf@5RaNC6H0aJW<2V67a6\X<#F7XDXW
UK<&G,Ff:X>UH?J^]D[OF@&f?K-Ad;=-YWc?]7E@_UCWM5^^N2eY#:;eT>@f_@;#
]bQ1L4<.S-@1@=2MUVJEc26-NXIL8\J\L=:5>-^#e_>O?M)ZG<&K+Pf=?T=X#<cg
&L:g9c16bfZ^M3UP>7_2g0)?A,\E^6HSUQ1][4Y-3\]27-KAB4+27>cC?K5QU7:J
Tf&(E/Z=H^7F-8dBF@@,IeJgPEX7;OdYS3+Q[,YcJ8Y#Of()_aT.GUAXd;WBDZ32
Og3d>\OMcgUX18?^J]0=L()Q38A4WfT<H8V:&3#;13ebNQg=X2W/<HD9#+G6M,af
g4<Q/K+Z-@H&R]7Tge&RW+G5+YR8IbLS^ZWGHS7,f\113;&C]OTfB-Gf\-A^B>.d
UNQ7@K,d&Yf#-HV)0Sg3FRO3KVG)NF^=(5[fM_R_Kgcg@J+;47I-\aW-UeLF>2A@
P:N_>HKHI6)b>:0Z8Oc07E9Re1Z-_JG.I;b[_U7U4X@6IB=X[++15DMJ4V[@=O0Y
#;T4V@V<@c:&<9]3UV\4)+33G5D>ea.Ge3J>f.=d9=1c6<Q.@ROU+(bJ,06Xd.?V
:82B0MH<D5.W1_L=C+SAa[U?K1_,;b/4#__C<D#W@N)/^<_Z[8Sb]d=T>9PMSY8@
60T)+HZd/WM>bH_WQ1;IW6a:WHHK>DX#XVPA_[HK1C<<1=g<b>+J_&V-_S=e\&_5
<S1Q^eYM<a:JV0?;7C6^7IL+MTb2aZCd]LT7KO>9^;.KXL)S446JQAc:UE9Y-cD-
C=+4.==A[T0B9]:E?NIM31NScE>QJXCURDT:T;S42O/QfJaM>,NA@=;GA+S/GXTc
HJO[c5[5S9Ab(;6OX/Z@(<T5=^gg9.G;;8I]OW.f^/5I:1b#.Ae?]_P;b\.V;GDR
58QgB/&+?MK92fcLUO[(PE,\<QZ-B2BVVLQe87V.9^<2S2SG-.67ec@dA)Z=0Y8#
c]dfVEfH#Pe7,L3bHSdP[2>,OPTL=._f]4NRfHAMaP+-?:3?dQ5Z,ITZ#DYAL.Mb
_[&^G7B.KJFZBD=_c0=SXUJP3(A;R3\M4>[/0c-8U;T_G06,7U&.RG\84_EXW]F8
0=0IJBaWTFY4:<QZ#;K:+NDPW\O,JDW/5a;.?:F)FR#<g79;^/=GYO<R/PBd66.E
:MW@M[^^@^L/X/L1W(4,CL9#RG2CR.DFg1BRFP;_UWDQ^F271f]SK)85?#aI88@#
Za-3Ff48Ve]7eER+MDcK<LA]MR&65;T2#VK1S4.7I5X.e.0PCS]P34Y6JfbA=0Oe
0]0\F([aZ=-XZBYR,7+bbPY\92GVa\.A<fe&f,PG6SIA6OMT0666aQ4OI)(M(#KN
:4X_1e<#c\59T>@>>BSB>:=O8\YbX5(MgUX[H\fI^R85L74b_@,&H<<_@?\SDbD;
#FW(2S>PacRW=IH;dQ@3=e;aeR]=LC78,Z<dAg@(dS;]5BXMIIZ?_ZPXS-=.?Q7D
:=X?2\Z2(5Ke)):B^+K;A64e;/fT?44.a3YG.bc(gHWF;/_#[FGUWO\Pe;KJ-5;:
>[bL?#O4OHYJGSgdQ[362I-OUD0.1)6[dRV@5^a2I/7Y)FWR2<H+2#=-1G^dR,\B
(WLcJ#3-JXe@B6YfZM&P,CM&II?E?I#9EN&,]cb[dG)8\H\N1&)Wa/]+&@LB6#4a
==9&_Z<1U4<?@Ib+U+).0:Y;]ffcWAe]T];]:QO<\R[dL?f.e/<V+4-)(]:)41#1
3b/eFGWO0eO=)8C8;,4b]<ZTD#U.GBX;GLX^@Yd=WY,J0_?T^Wb9Ta[Ke=YD8EC>
\@fdOK>aW,6bZ<T3e8]]W-(J+7g;JF(66Gf#aBPfBD0cATEZ;;=9^38P-9XXeS>?
&aO--E@Pc(M_7gG]2-Y@927P;dI+aJ99N4M2T(Y3675ZdJ4?Y\@[^/A5=bGI8=KF
WHI)HLA7&^NEA,S1J5UCERbb8;RHMM8NY8d885B0^7&HKTTS\2eP,B=TcV=d&IXY
;(J\aQKRYZ;+K9WV&_a8[&JU@@PGcC1KNd_8C;NN/:(_@#ZDSQ\@13R[83_^c0cf
17NY_8^;47R(.WLc4?Xb8GgR;;2RTD16>;5Y7-U1U=)D?\#>fC:_W1b;<-TR^f#X
<gTT[>;GJPZ/LH/(VS_]NOW\Z.b]S78Ha0#BaV9CO.B5a5Rb\^>:8EC?L5)R+RRY
9N&,RKR6a7.]#TDg>X:Pf/g:V5a6&]\CfW&W@?LUI:V<g,g,/7Q5NWMGNeMf]Eef
&<J22,d)BP[Eb=CL&G.Q);K,NFTY?8)S;[OA(Q]BRCSHM\^fRBA>JCPG(+[dEfNA
<D)9,U#:>:=][SGQNfB-fIG:32Z@bFf<F2P6]WWQH9/<a6KLHSP(>FE:a>cJL;_V
2Of,WKEKSX?#H.Y5,;3DDS6Z[Y=:W&E3TgNc85FYKgV_8a\,B@1BG_FOD3>Bc>db
A+JJ.5R-GD>[#B_EbI&=aY9L?ZHg<50B-5RgC1?bRYLGg0.4gefIa9RN.ECY@^CH
=7_N:OZ^:]?U&@.Ee>OT^<1;3N^Zf:=:cWCLeJ_9(([GXa6I:Q_Q4)R6^Zg,I3Fa
/#AYXM_6ae79TKB8b/V9]4e;^6>-6FdJ<L(S],RF-4&8BEQNZc^>TAB+A&96KTS8
?FBOg+_^d3=C:\cM_a2(5+W4F<Q&UQVIF)KJ\:UZD//T]K<HPUOB25X=\b]ZeA71
e^6c4V5XfbG_T<1_L2T^CW65G>ARU<O)WIQ\(@.:G=aa161I?7^g5-FN<?/SC^,5
,_+_,7^;P0H=0OU#bD+?AUb<;+;E4Bf4J.3c]0G</#cbY2<\1Ga:Q\gLMM4eDJ8F
VV]M>@#,J8+3W3U.eQG1IY1@K[RB:AXeNVe[3ZU7F)&]2\Y;>:g#S-&cd&J+<C(A
7O8]<V.<\#HIDC9A0Te=FM.PX.90UAO(LH6OE/#K.)_3^B;)&6KI>70.@YKT8>UB
I#JW2AFWaAe/W0;TU9)Y59f^441P(4DED>O,4)O,FCE<TaQO11.JTDM2<YKIQQNZ
,:YdgO8V1gfGWMX7\^M)>P?QU>LM&e3MV\RJ?^RKfMVaLV_KB8G?NL?.KL65P54&
JHKM/B+4GDfRU5/Z9\^GFQ43_/+&Q68gL-aA[Y0J9:40#PMM3QXL_.2eZ.[G2+PQ
>Y+=/5S;3#33+,Z>UD7A4gZHJCFG_KUV@W0W#8eb&L3],9b.1G6-aQ5B.NDb,<+:
DK::AYge;1c^Z6d,C^6d;VF]>AWJV5&#5YQ/E0-eQLVdIW?e]^BX+:f->@L=DU:5
GL0=IM_7[=E\FRW0UA-Y?b?cFeFdQb<X:@HQ^;QOQfUf=U@N>0XbJQPZ3e>Y1CI)
&_4P(]\C@COTARO4EXV--aSGDUO[F?-KCIQaT,d-&96TV/GNAfS2QD+V+aeD<^+(
P9ff,\A@8P?ES&MI0ZZS;7KYLQg.<;&\1K2dGI#\Cff0FCA@KY9fd:?KKRS5<&8W
#E/SO+--JP?U8>+O2aIY>Re_2^E929(RK[Q#Lc#OU.NP;fSNLdM;b#gL(\C[+4_4
ND?L[8>H5?g\,VE/A-;+8J9:F<.+bFDaQ@:e2/GFG8<@He<2(VXSG8Xf18SS8.4D
0:K>K^(._a3dd(]X?I>6&Z)E&MI:<K;]B?G#3(34&GaeIC9P0JfM0]JM87&J7@-<
OeaBTU8Sc\JZI.A(g3-T)De<^(f(T45P)W[#S._ZCP>).:9HcEW\eeC[IP&>eWT\
?MR,9Y@0eL/6Cd7:,N-(-I21_^+HK@_B[BT5ES.#:4.D):_&J--].QDS#=R\>I8L
>Y([6Pd_)C1SN\+KY25\__)_\2D[&UMeROZ#[GSg+-O@3eM14@P?/b\2S)0ZV-EW
-W@61&K>/Ng:^88f2E3/(ZTXcaU#A@7X)4A_bY8c8SYQJZ2Z/)9QSUF8UCQ=_(6a
C&@]FRIQZ(:af:.f0]bCO:6R(K<GQ+:SGF4:ZS+;PYO>3HfGVE8BWK^a#9;OfVY[
c>BbJRT3Ub\G&].:FT?f9cW[?[HHPE0SJH7c0U\?KS+RE=&Q_U)2EU&gY;(.(&2F
9I3)</6C]fQ,D\2M_T>/+T,79+g5KK#Y#g\\T\dQEL+07Y7EVaR1Mf9)9T67RBTH
<WTGbbBca(_@V,2-5WKTHEff3QJ1HTK32[(WPg=Y6(6aF?:0E2]E6=4/L_XHX2&R
_4#,>L_<NOVS:[>3aR]FZL])KYP/&c8@+E:8@cXZE5\EC:)3^X<(c#T8GXG4)R=+
<MH8?XbeLb15:e;UPMH>#cW8S&V,b;G)IF?dI&9BVKG.8[(XK>MA82MOO:1+#FV+
122cJ<d\7.ed8Ng?EA4Y^E?BM>Ae;<MMN?]R-V\>)E9N8ORNM(3D53:ITB<7/d=_
+60MPH@7>4_QT81NXAK;OZ@]E24Oa>#K8,\=NLbP-8a>Z:3@G21/_B.1^;L@89SC
2;S(FWV^@#&#?H#N1USA+\A)G#AB>J,)0a8@gb\=Fc>1P1f/DM5,bF,QID\+Q2[d
g)P>+;aD8_Q9_5>eaKLcCK]WT676a;.)S&D>0F<Z0:SK6DOUQ3##Eg3E3T=AE1bF
-[\(H@VQ-[/;B<Sa&1+0.c>NHUKJ7?K)Jbb_T/dd0P:fX;4XUHE>d.<@Z^0))Mf&
B^UaF;2d4OdT7PgAf55e;ELU51/I^.]5E=5L9]8;fB(^?C)M+Q<3IGI-W?ZL=b0,
KB2UQTVe017@4:LI/1E#XEae[TAQQ@LQ4YG(=7-Aa39S#&I=\VCCb0Jb+Q\1(gfE
7\T0g3DRJa2>M8BWU?,EK20QP9/XH90Mc=4ad\JAOf4?-\I1C^O)5DPT=RKXZ0;C
aS+B],N;JMZAF2395ZQX9V5NT<\#a62=b4&PdLNHDK&_V54BQ,8Zbf\WR&/f:KO;
eg-)eIg;)C7[Q&>RG#6^#\#<5g->=f]>/JX]W._Q)24<M,CQ352&V96aUD=-]H,Z
#-eK^c=b_T;a?O(QY0-f9;X\f<V_N)-A&@EbY;Z,-bT_(6F=8HB.MX(KfROC0L64
S&1f?7ZHL_8D]1aB\S-W_:N4QMDLY[e:?7C@.9Q:/E;@&VG8DY.UI=H7g^@Wf(\)
=Y)75f&BKcWVKWV2#fdA8-+gIF2J6eALL/b?ZTIcXN&f.\_9a0_<d8)UMFcZGX:?
CMJR6fH]K[WZ\#ELa,RTWR1,C:J3PeJS=CSL;g1Z1PAd4=e0S?\?5U@Ed)>a&=)[
25P@.L\<VSCA\:ODMS\XH]<F1I<bD-M>S46]2_I1e^L3[6),#[VdIHF[^,4(E83d
7_QH1G2&DF)@L&)>M.GD-4;^G_C;A^]V8,Ua:8/IP8A1&&X.3@[PZE);a^e/Rb<)
46\8[)__HP(cdf_39U:-3fSa)@cgC1P74LT&09?1396IT4<.:b[.XLf9E((<fg6:
BGf/9X>N0c9W00)Z/U6]A,Y094Z,&KS4X[IY(EIA=g-(\>U2AH/#C=8Y?fFMY[Z&
CGLI5?&?O8Q@(C@GSMecCTM8P75Q-S6_G>,4@65D(3PQ\1L5?F_1eA22e:@A8J=7
R:89=a)bP3D[N1Q@W(;e@-N<[6WDV7F.8R\C?]:I[H)g&)HL[1Q@e,OH-9cXcBe0
?()RFD@_@/d2W7(8+.>C84JD6NFJ=T(HZRFA86]F4P_QRY-5?;gN0=3dUN,UL.?O
V0dVZIcc[K@RdQ<IeE:Y=I5SWC63Ndc@D]eZE(I-E=+)e?1@N\cg1-5/K7,.@O=/
2>77Q)F.U799([bEg2bXb0ZXd8#K+.J@gL+N6Yb4DHG)[_gSfMYN3G3aHW9;M@-c
WK,+c=1^a3Tea66:-gB9,H]Oa2DMO#EHXK2U(LDXfIeTC7#HRCY+Y^_YaJ[P2e+P
O3<>AP/\7BS\<A/gXb_[<,P_5.eL]eef,6]3;Oa8+M7cS5<S#IL;B\&WZ77-R\H/
IZ50+(BJ0#GV-3?;[.CIc+.&Ha5UX9;]X&4@.4SC(BI.PL+5/L8+C>cM16gJ;M__
f=1J3N6f21J.&BBY)/P)?bD[354733TUOLa3@_EU#JNcgdf4&Yc7:L^JZ[6a-M#@
[g]G->fSP@#<ePA7(g.2Jg+IZG&<W[PK0d?&_MVV6FdEE<-1;,73Y(HBdC-T/2?@
]Q[dJQXH62<B8JQ+:Jf()cbG-<b>A8#T/)05#-.g>+11&T#cW\Y.5K>X;M\_DT1A
CN?P=JX52E@)/<IJe)68>C91TAOL@Y@I;0&\BSQ34J^SL5dfY+FI[03e@?K<X4/2
/X)WWDJ9TG0:g7WJdOTaU?S]TYVQN(c,CMTC2-,?Q=GQCYULe5O)eWT0a2:4>+b:
\[?^7d6#_eDL/+J/:XUHgJQKF?+_)fKFX/BVO=6:?cMKD_P]N^UKS^,C;<4F_\GP
EFBe^\HTcbA1PabF(6-;82Y@J+RH&[UP;8]+\K&Da5ND-O^MY>DR^M]UaWZ,cEXf
RU=M(0X-;<I6Q[aYO915HN.E2S-R_^JLW<ZfQ^,Kf],SP3Fd-&;(e6Oe5<U4N-HG
YffH#7LIFC7+@d@4DQe7AeFHOf]XQCd&96+OcK/?YFHLGV[bK9Yd58FSCZ7_I>K@
4<),fQC\Q8-f\?1d@ZK5^K#O(>0gE/;,/\Q7\P[./&^J<N6e@,L0ZE:YcC@A]f20
ONEP@f_E?H(VeR&Z&?DT>O-ZS&M18,(-ABBZ70a&f+57VI[1J-:5IQ6dHGNP8^L@
8S)6L+&D,,WU[C)0XA48W.+,g)KJ<FZ1@MeUW@(D<)FQ:gNJD.]-Wb++f/,UVGGF
[_fF]MFB6>2Q9=1X<B1260TUC5G?(b)5&Fd/1[26S:+.C>Be7B#OL+.\O\(d58A3
DgDA_VCKT=+[1E?,=.<HM)88A]8+QZf?=PPN596H,6?V]+@X;\7G]D\cYSaJD9QZ
NI-AY(I[Oc-dPU;6e1L3#TCF.2-CaIB=3VX;.Z?dM0@I@c,Q^:DAAF7aU43V4b\d
A>a12AI710:\[gWE1V#WZf&9U&6V:@V49KA+>1>(?OcC9aORBC8MIVfYZ=BbAJR7
)V?9?If\\GKT;[f=K?Yg\YTXKA2\+[4OUD98PgXZd6QGfLW8?]Hbe+I,98]V&9:5
).<M;9&NLYGd.@XZ,UT[,.:Wd_0ZMY#J7M\HTE[>\g)KRE3B=]\[YePf]bF.7dK0
V]ef<6Z-C#I@]SO4YgPg#MZGRY/a?:>?]_>-;1b7MQ];^K@g.O.7NJWZ8@91&,>B
GL47](+>W1F7_HS0G5F->L)WV1QPC6S00R2BXE1F433HIdQYY.4CWQZ^.PVNG7D8
de[3dcEF3)JM7<aTM]M@ZY8YNTeTS19G08gc_O7_OK;d,.GARZ=66:)&d^D[PZd<
G+/&A^[24ZYL)8fK?#_8VJN0H?BM0;Z_C?F0=Q:^9gMS&#;^VGKK>+I(+BS7,YAM
ZfZ=7=XdJ4H,VH/4fabC^VY>2_M1;PXcR>Z^B&KNf2BfKa[e7da0S7RdBE]X)R+J
Y:#4G_;ET1I(FW5;62f1Q7F6_4Tb-U>U6JM=#&GMMVG3MgQ^NWEX_b^^45@061SC
Q,Dd>S&B12XWV&(4M4K?Cg^]DT^N4>SQc.4#\e.gb&?BfK6(&YeWQ)<8\Q#IYH^Y
NDHY,54J5NJSE>QQEK5aO0ZYF)-Vg&_3ID-HOfc5VC4BMVY:9L;(#;dCQfOJ379/
f,>.T)@S.e)[L\C+G^5FF4(FOWUMGCHNQ^Hg^6WbSA>=Q_ca56\;5BJA\5/9Va8b
.FL=(NK4WB+0=(<4eC_>;6L7#C_=9LF34638Jc\cPeD;,TRTAC&C6NZ+58;P1M@5
?B3Z(=.5HM]5^<X=PD]eR^WQ=P^^DYA9f;HE@)3--T5^6C,c^CW[JD4)3B4F5?Z5
R4K4@78[?AK_eDeQ7?g57eQ_O.P7EQEE+;Vb<LXeSc1>E:?bbOMB]afRUUZZZNO:
^O+E<[JCeP-3g5a.UKC)Q82Y9[3-Hba,QUcFOFWGbNcN/LX]:@Q[LJW^+M\^)@Oa
XOL^.g/\beQEAQ[:+X80_Xea@;LOJdKgC.J&.NQFbMS5OGY_ccRI;?+)EdW=(_L#
Y6^)GMF5H+e9]G-HZL\Q3AL-#LW:>P@<C3LP2^@<25I155&43KM#X2RT)SFR;#TT
1a#[XX,/XE;5UR/=++HVQHG820NK>-&-Y15G7VPS.Q_c+?YXaPW+(#J,#Y736[g,
<6>TUfZT3dY/.#JAQ[68=&2<_.0eDDJ,dWRT0d@GVH+9][;Lb>3#07:CU#^S)I+]
TO>;@/=TP,F4CddWAA5-T[P+=U(\K2XfNTIOJO1Y>KEZWc[UCNQNaY^gL988BSYR
QVYAPGE,^BP^^^^YcMOYS/6cS9R:C^&?#1_Rg3L2/K^#SVU9=FI^_Q&3d&@<13P@
eJgUVOa]0:/G#)I-.e#BXD16)gT,Bc2-H#E\/(F\IM_7/44b&I.9FK(2T_)MbI<H
</P_OG2a0K0-Q_b@CAM+PC3]Q@)Ec\G(_?H&Gb;S<T430X<[1CKS&-O9+AA?MAGV
_KAAd[gF.6C),;[OLKY@PD<I(NTQ,Ce8X_bI/B<0ZPD:TC:Z,C19>OM?D\I0]3#L
cC):SAY.Y8GJ;8TfF[+:73/P)JNW(194\3PN4JWFd,DT:^-bM;dC#1/+S&\-1VPa
Z?^GETI(7Gb3;WF9L5@TJ&H0Z(XW7M-RW.+KC+VD8I0AdKAJ57(E8;]U)N+/F1_Z
;[VI[]4<PeWTOI^\._&,9-ZYN)4S&PM7G,#YRCa0M/AV?Z(286;LY(CC,RA7)cH(
W.59ZKZZ.;TW77f\-JX@M/4gSO)0XER-M.OD&a(L^SP:;ag)._^1/UX\SB4(bHde
PAd9_CKPPT0(UM@8M8X9g\MdU8)7EE/Gb2c-e@RTc+cBIe@S-V[A)M=)11+PdE(/
aEB0ZF+e,eKE_P#Pb-Z+9Z@+=(\=#IZU51EIN(DD-79b.&D4_I;DZZE+TF,QI;5H
DUFUD(]>D(-fFQfc-#GQDD_KO[6bW)9=L&+2E<TbW-,.6XPC[4^:PI46V13P5]?=
KT)LAXfaL02R-NB7^G=EeaD[8g_R6&5,OZF,g5.YKYNIged;=0G]CeUA1a]We->5
:S<XaKPLFYUTX<P@P0<G(7IXF/W)agD(bQ1\JG8bO&;#<YI&dA_^YVZ1gUabTH9:
dURC@[5Z9S4&8,PGW_SSZA/EBK1#V95&/-FIM[WXR<e:QPAQCbVd1FN2G6G,.?:6
&,846&:3F[WQ+5N0dd@]ZY)6;#e6V:V[R8R9]+/gU2FSgW)fDQFE\Q[=,JJHEf3J
<aVY3M/VRT-VNX,Z;A21Q9(9WWT[Y0<Mc]UQ7)JeCC261dP.6C<23_B0;1[RM-&&
JAAIU_JK+CE@[Y-,7.&QISV9@[D;BBRNP2Q<O8BL9SQV#@=O+#PdbT;R=Y0R9;a9
g+3,J&,GTgbWe_0W(f<ON;4f;BMN?IA=D3X;=eO;[(a=WD2=(AUNP@(37(1\=OJI
_-M[^)&3(^PG25-@[ODA7W[GVF^)LW8.KHZbE-Of.N;1,e8Z49_TD78b403d9:_a
#H&gZQIFM6S[bL8QaUIZ=_B((QBP9Z.gR2=XaOC4L/>FLF.\L-M=\I9A]W7GdfCc
-JO[3D;EWVEDIO0A3:NNe8PW_\CAS8f(3Re#KYF--c\(@<I.;5\IJMdcB93OOQeN
Q_5Lg_-BHQd:LCVLOCa_ffNF=-c<G1KcWJG#7D&:6G<0W184CW&7PDT.:B-5:3fT
aP/,d7#OS_+PR[eRQ[?-G=&F:a(+f##41e(83-P+Y?d[c,8S6SdUGC=P#f;DJH7e
OR/@5eTX-^:bMb;Lf@=;e70N)bK/M()c3ZJ7+3fJ#YF@5)N)T+XVAVD]XT<7O6eF
=Y34DN1dMgCdA.YcI:a?2cK)(;;b_)[Oga5P6ePBUXMJbb5W.1Ud,AGQU24YM7LU
^-5(]XIKT0T6Nc]HeRE?fU?1F7JaGbd:B=MXbUOa&QKK,R<W2\8?..9@M5-WD&0(
aHg^:O3@>#Y)/26(gKV(&+[EK]JP[)[--F::@dP^BCEAegSW0HCN#cd>MZ7A^;D/
=2^a/#,.-WIJ:,(QaE5NU/_\g:MMR.+aKF.6J/:g+PfV:dK6gXc:J.b1e9PYC73V
3ffgA:)6UO_da^Jd=Qg;Z/Mf6U4;8W[S=/WD2JLa>@eZ@CC+]ec/Z5(DKV[5bMU3
H))6)BHNH:9PBa,,\0(6ELW&gK(aUX(J-M.F@K2\FW3XEMYeaD&,g;W(f0]L^M9O
Ug38@@DR=LL.0;F([;=E#-+a^,V8&[)U+4S+5/]3c+X=MH7)XT)eLa:c7P&@LD)d
+45cTbU2)-R8ePS,3,Z#NUYFDCLSO>;-9X#N75BGRdVCF4^^caE<H<DX?2a<>IK9
]gg=)5_UW6fB=ZEM3eZ3XOa?S2ZeRg)[TWa4aQW<@;>Q&W?OJd9Z[DJLI4;&I62:
);JHK?3G-e&Yc?-7ebV#+#?6VB]G-1UQ4H>1<5a0UgP]]>(D=?>&5NE@(_g&.E@O
N#C+&I/4]bR:&BLZIZ6@LKeH9C0LOf_:+:eJZ?3[9CEW[BReARH-7E8+SW[c3RX]
[10TS35eN6FAP6:L[Z+Q&)^-_C9K[(CMg9JXT(;aK1(I?_VDNZN3MLSJ<N/5E068
L1YfGea\bBZA1;;,36YUV6V];d56H2B::BJC4@5-D<_.]bJe.,Q/I3N>-DAWAa+Y
=MHA_^a)TW\I#1210,^>:/U^5]_c@OX8O5.fLgWH=]YO1JeS/c#];?,GD^df>4O&
BTRT@T:f3E<:L^FC?3UAg0E1bX,8PD2ONd)I[.&EKO.V>-dV48:TAU@OF,3Bf3;c
a+.4FF5A=U4&,OfVH@IDE?b8Q+INg;?]R3OSZWE;c^U39I&5c]UNcTNV[UP:4ZG/
J65Q;X.gBVN7&BEG9K1U8@SUFb_LZT\>7NPFdG//&K]E^1-K>TJ0VR)_#PJNO/Q+
(4G7&@W.eFVfb>J8UgVER.@9K2^aV(7Q=_;gC9^b5&=FAJKJ>M;bd=.0:N,R&0<T
@ba?GK5L4I1P2=MRbZb+adBZ&c3QJ\</fb>/WY<bD\0/4^E2:<(eVY#_0[9eLY7^
1H5>V\CV</^;bb;74>+T]@+L9BKIE+KU>@8DJLL[(GG7B5Z<2d#-)e-1[:^E-6N^
V\:LW#fNVg210^PEH]ObMTeX]P036A[=+c9H5#OI#:;1AP-_&RJb^TYZ:c^WP^9+
T,KZM?>L4;F3\3,/@dNE6c(TVS/a:1&&ONHdLA(<4a.gCL2F1,a)[Ee0WAEGA0^,
&@2HR<#QJ7)7Z-@/Ab2IKbSc@2_bCfY,1@3J)EHFH290f.>aYTB7.Z;\cfX^KHB]
3.S.#R##MI;gd&<U+3e>UbDT?.CNLX#8P4c4(/VcN/7\/IaU)7]>]R&WE<WF.Oa;
3V<G#X&KE_7ZZ/5\G&I1^IEE:GG1:JZ3,TYDRN5YK0V](#[V]UO5R3c5UOFURg<9
O[f:ES]PH^9AJVR_LTE2VNE<B0X3/[(BK^R]T4Y>^aSQ>dZPdQW]^Y<HWZ>J#7RZ
BT.NLKdQ7]=b(2PCSI&/Y>6O0+[5G08+?Dbc(3dM39YdNH4EU8D\HK#GIF_?J37Q
_G[-EHRbD=;4:SR:&6S5S(Nd#0b12g@@AI2:N__2_Y0NfRK)35)/?J)>7b<b[Y;N
(<XP=-b(W=ceZ/BXQ@U:ag11#2Kf#[T6DEGF:PP<>bHbfQHGB:#_LaQU:[b(aMbd
Z^c/OS9&2>>5b#&ZCF\<BTHH2+O(2f2,9Pba<>\4H>+]^(IWS&=+QAKI0/.+4_WE
1&#\1\DTf<b1M7QZa3K;BQZ;6^[N;L@cB(fJe82?1BUONbcB@1ZLJDFI@\^2W(&;
IB&@0-[>^O.[,#T/](ZfA<C)cX;\I)TX?SUbXZN#d+?/(K+,@LX[MRHaKYMB24J.
EDEPgQ(>99^33aGN-0[Q<cKdb^?H@Weg3DS)YY]e4MTF003;a/ZE>M>[V<UJZW8a
IaG_3)gcQ]8(I[aEZ[-HeLMJ8:2D[eO_7,/)R^(f21^Ce](S=>2.L8]0Kf.K44Z6
[:I\MTWJ^S>:]<:#YT<E]AbOGfGF./XPU\Y?EU&?,D<:1[2C&&T,?E.L.MS12JK^
WY[;[77;0_1+(-XMOOJcC9D5,cI6+#eb_VE;B6N/WP-+=La2,^84eX>HR9RL-afM
O5]>-Z\Lb5^6fM<e]YG#K2TV;#>a[X;8<NM<T+^JLS+W&2L.9O0c?G/P\,)04\_2
B;LA/H.cK>LU<-EY\RG^A2&055+B\-Acc[V,EOMOITK/50\VKQ)9/Pb)USUeP?OY
7#^C-1f+ZVIL&J3I/fWB(3].7ebaLLEd\0cJc(6QddK])8]K6\=4J1L/KNaaQ<F-
=AKQ+P^M;EB5c8H[f:a8>aD=LE/,S_79TdZ/0ZUQN&)A#V[a@I.7F)X7<[Xg9JgI
0Y;.UO1[N2QV2FgV#,UMcZLMQBa@QPJP4H8OU1&adBTOR5a=8M)6:<4=Y](QaF(d
=4Zf;?179OU:ObRQ@TU\\GX?(OVLC3Q\9_9>Q()Y\Cc0Nf;+29d<,+ERfDXDJYMd
W,\WScVPX1=[e=JBR3J-MUgK^?:+SfLP2I)MfgP/ANFaUg+cSH--cYTDC#?5Jb8,
3LD3-K23::>&N-\#JfZ=7F5[HTeK#V:/?9BZ82#M)FIa):7KQec1W.fJ2(&>TSSP
d1YHgEJYZeEE/a1UMg(REdS@TA3K_Y]KG/2O?4;AG@L(_g/V0Q=P-EM)8KEb-.PA
,UV93;Dg2H@??LVVcad<4W:dK#OW2aBZ+Y;YAMX6HY/G\:#>F\:>CHLO3GIIb0T&
U;Ff5aWMaJT:f.1ZU5&W.8@c1e]7]-@SZWU)=GP9bSbc_TX4-[3d2SK^QL55MM32
]/IC^TW]II_(+E@HD25ZFRB+ee,(eXE<738K71,PW(8=XI(:4RVAc4PF@/>O;8Z/
XR\@DX.,e.L^TBQ4V=G4N(145TD0SIUT#XE;egS;QUHE9]#&>EGL0CA99GA@Wdbe
V9K10N&3,e+E6HW^NY;>A:@,7c+7+\NM+(S6fL6993?O45ZTJPbJOW3Y=4DXZW-(
1ZZUV57^fW9d3M9#UF70/\@5JW83E>V]J-Z@GG)]I;8L_A8NR-DPV+M^-FLAU<[#
agM8#;\U0V/[X9O-(WY<IJ1F#LQ4T>FdE:f5C8&HJdM[4G7:[E(;aR@8&DPM1YT0
P2PS,M2<T>QMF=bBfG^\3.8((-7EJCFF#+-aI<I;d5?-eXK,Z:5P1..>EbEBT]7c
5CF80,ag3S9&E7>[)^3g(/EM8W.0D[5\QUVbfg[>e--0(6M.X(D89gV9H@Y>GQTf
OWa/P75)2eRddM.W3:MZ36=[.N[=gEWZ6KTO1fHT^\CBBC-fRP\bT\M>1)DV57/F
EV+dXI+A-^g&bG#)We6T8U1J;@=Q8Wb/=-WR\@cB9)b)N\?6S3-<9HXN?AS/\_M4
fFa-fb4VW-YR;2_(M3:Te_X\\&\Q/?\/(?Y1ZCPYdB+Xgf)X)M9W+YNR+BN+TCSE
[)<67Y.GR7V+[,;a]VDG=STNXMA1,Q5130=b-:23FUA>V3>#Qb?5;V[RSRFge(X^
Ic77;AK2>[IC,3[YO]<19@W>T9(?HY\?Cg<)1gCS0(-VeKJ[?NaeT31Y;NTN4B.e
eF^W/)RBQ-7CZd/&:;Wf0aB<T/6Nb\\HZN/L@Z;GBU.Yf1L?7O]NKE>Z,bEULN\I
;@:1;Y;)[E>=?L-HfBD)H5Q)Vb:[EV:);M8&,Y;2)6I/A&)AI>2#^d.=A4\<1\2g
2g2;cd]>05U+H0(&+S:^]<U5B-S=#?9cDeWY#5V-?L/Y6NJbf0d4]OO5P<E.TPBE
20b\I?Q:@&Bf91IRYeFWWX[@RVV[SdT2=&bIMd=1?33JNG/V,U,B8a@9O.L\((]9
[,D5/c;2@PH9,N;DP^dD+ReN.Z#OY_)VVOc&8W1&d(5^fgNTSVd]+7]&e:a(SS&S
,I:^W:b)gIdYGAB@^IDBC=C-O@[WMQRJH[=P]65DgUf._RFM[H_44-/.?9I+?224
T5d#5C1&LC#T7J1E31?Y#T@#A=UDa9_-+_Y/d:&/aE4dAA=b[^N6,,.e9U).=045
@40)63J8g5Pa8;;gaYTaA+[g9#,6>,?N\cE=E?YI0)SfY@9A1&5b3fX-U&)0JGSD
/A<A=QKePYM<CL)UI,<\ZTV7Ha9#@YJTPBS_=cd^f-5Z0NNCUHe3R?F@JB(>&cZT
L-;5,8&/G1A\O_YRg:f:e97RE<Cd0b>QaV.76ATOS]XF],1RL:Ia31NY)QJN9&Q0
ET:AJ:4TK;K-I/:\[7N-,&<UcW\)E<#Se=C1<E4&@.;dJ4TeNB7dFNOS^N=Y^DS^
-T#ac5YLU@U8JcYd=P[4-.OP[9T00\3a2d_^\S]T&PP.G&-5M<\Fdea:NWO.+5&[
?-?.>Z&VeNZM@]?UQg589[J<UR9Q0&d@(.]M5D_2GT9Ob:#(+B8F2DTQ_Y:63SS^
VW7,5GZaDD^EE_afQba(=>Oc/K2M-HO2XHB=,3,VX:Y]9//\)7QR0H^Ff2XX\<bL
#Le):N7b4I,3N)XGRL8+:8]_]J99,H=8:bAU65]KDa4gDUENC;8>J9d]#Sb;F=ME
)[dV4e/>^<Mb9>W5[-8NG;4\[,cM_BWWP\<-PgF58-(S]2J\f\:DK^3>J^cH\9NO
/[DF,&#I\+/X4;D](Q6]1]^>c9H=bU8-+AaF.ACNTC=^2/,B9QaeEA(eHK>@64-F
H\I^N+5<#;W6cMFS2dg^;_GSe3S_LDf5)-X@YcG#6DZF_.QORJ87)eDR.KTb/,LI
)5I@;,dS#@31(-=GGIAb0QBN#MfcICXP][<T2\^_+A00eL>O#A-J/18,e\Ma,GDc
O<]=6^IDA0^LQJVCc/QeTDe.:U_Da#PMTf9O&bB6Q)dRIMHfOYL>#YQ\?>MDV5dL
D::7>#N&>:B(+B11Se]4R;N.KT9O73P]:abG[?MP[Y7HgZ:Z^/+LG+]7:1-=8J&>
9^TCL/]ADfcW=UbCDf?(ZeNWV7NN255eG.KFL=BTeRdfKf,VZ-&\HbgZb2F_>f3F
1KX9_\E<&_XA&e/Lb7/V45C7e,ZMEeCJTJL7@Z-ZAO5+\3]RRL4<RR+-=PNAW#ME
T;.:@3&&b/,E2eXPA5>&3./]0CRUVZ;&A/-e)RaOcf0a?3:Y)Q4TKME==a7AdV^;
QMJY&1<(c6C(92b?Q-E9RBY;7=\e]eGc<<846BZ96Ef94\4\4()G:aa37e#/<O4,
=5-2]8.ULgVKU(&#F:7.X/T:?5RARdI3dJaP^W-)CADA<9a93+CgA^TT^\PF.D?K
YgT+P98^FQ]Z]g5g4?B>a]\S(-We[0-QFLN(^=PJ7B@CJH_3TEKb80cY@?O;gQ]B
d-gE>[2WL-WK5@@DOUY/b3cX7FNI;DYOAge=BS3-O,8bc#S#UH<6W[aI06fba0TT
)eA^b,8?TRGY&bA^MYbG<#V8:)g/8RTK#_[Y#VRcDG6Oa#c@N+=..)&K\U>_N-BB
(?GeDU=Z;^c:=S8K/f3Q3>\FC:7SE/W<A___e5[\KOc(N9#B)VS0;B7RU@g@,GSA
TW?#]e;>ddFTL>f_b>A?6E:7JF)MLI.)]9XSdec-P==M]GK4<aIAc_FRRN[RO.aB
>RaR@Y\LT^ELfI)3)-T7D_<J_ZF]IQH[UW>D;34L;)K)^Md/[7ge]J-MG\+@H\cb
V#;DK4dJIN?&gFT)CfO5#3[8T[^g[B4\@L#Q#M]7b&SM1U,X@R8+5&]E;<Q[8Jd)
gaW747UN^9Y\JG#)g;RHLd],^[d2^fHOB#_=HK@#V.<O6W59fR\^VIR)>Ad5W.):
c)JC_(S.KdJ>;Fb.T@bE:B]ec-;;gPW/..22R,eQ0f]Xe&&?R:e?dF@4UM^\;W6a
L.^<;bDb2T,Ve30LHc+HZSZJ[&5g:<>6(AM]ASUG@dO0[/?ZU:;ceMc@Q0SL0OSP
.S\3>CY2N,9Wg@9PM0:L>X\NXZ72[/ZLJ#@Y;N1G(2Z]NBHE]&)(?1,#Jf7/E-?@
\Jb#WJWO8,E9Zd+edSL#>Y2cCDOKW4+P8U5JgF^2[V1FIb2/Sg/=[9;>ET3UT@d:
S2O[e^MU6JC7=7(2]:1:-Z-dR=a=JYQT;4F>bEOL0)b)KOYbKX(9YCd7I1;9aA_1
eE_[Ycb\\0Z@/HM1F=K_&T4_]>DQ#C2BZ#,;]GM^8R7&+:FP2#EW.Q@C.=\,_:J6
DQ(1VgQ-46GL]0]DfUO&#<V1QR<[Nd/.b940)^T[9+()-cMN]Q:e[[,NgY\cfJW]
?Z4XZ(]BEd@&]eCW8>\=,;7<3U<)#&065X;g8cQ+Sgf<:LECABF/?4LN+9aW<Ob?
8(V+UZ6/Lg-a7/]DW&RW6=+VNEHV=Ob9<@381cb.Q^bAgd4^fR1cD&S]@KVTEE0(
3NTLN14Be?D.WK;WYN#ReD]N6DRIZTCIZ@d+2BB9_Z(NG8+X1?c[NE@_^^B,.4PZ
XDUF+/05S?gbC7WIIMRMF94A9eJKZF808W#M=)4b5TPT#A55dfD]9(V+X8>\BP1@
Z/AGb8]4VC.MDLPZff^N5,Kf@WI_^7g^2Xga788II@eDX/(_\fHY]65=Q]KG?Q]?
8?5bMe^1(-Y4P42-H]5gXYQ[A?KeHOfFDO;@AP[9NZ:gR]/Rd.H7eAN:O5J2[TWf
11+:7^3?S0cE21<78.E\+X7DTdGP?-?/.Q=1a@C>H&44NL1QO..L6\Jd;3CF5L[D
)U<aCC@0=3-E-9;f[7_]CI4?H=@9,H@(A>80T;5a=dP=^;e5f]D6NeB:K6MXU5,D
,Y4eH)e=,WDDZIVFHA8e#S+1B0-,.2-I6B<Pa/8=+>=Y/.^FOR/GIbDYA_[d0K9g
^5#GP6ZW->_#+[cKL1P5S;.SWOH^EU31MV7(Pf?]PQ;W)C4RLfI4Z4C4d6)fC[R+
<1^=7K(7QX@fAH@7I+/)_ELbY-c@dOR)C-?=?EOe:YAYC+S,b_[X7EP89-E/1>PE
@<7c=U[VMBg-8G)eK_\_+\]]4)8UMJ?)eTNd5PP-G75>:/-c4;LRXEcQX]8?WY;e
JXQ=^;?4/KLG4M73:,c+7_C_+J9N<?<_KEa2KR=6A90-O>7bF?YPg3E09RN\Me,]
XDOS=+5J##-C>eL^bD/=H#^1dT4b9>(1]QcLQ.YbK]SS&VOaLA\J/D/_bgG)b@T.
[1ZAP)gTQJOG1SPF^g+OXde/FY/LW]554-S&2O7&#fQ3cS@1OXUVTbK59=X.Oe(R
WTT?C)C[2Xe,VMK+>V>7-CCT9=EQ[A^;KL\YV,]Q1=<5BTaISR0XCAa0.ND7gOgB
9Da-e/BBPc?802AYD(_@1-N:[(L/60J?bY1[-IIC72RSEQ0MB4GdRO\BU)b@/:e=
R>N7B+(36MM]-d65M=P&bTJ,Ug=G70P3[Z3:[HXJ9ER5VV9^HMaCgK3WHY0?7DQg
PB<E[PeCKdZW.[]7#R&U11(2]9&Q?H43+DWfS0)E\4D;G[8M^1I2(GVY>B3#_[.?
[+2=(BWS_DW6A?/E?IcRIMR1=F7Tb+&2YZ^&F_R1Q\?Q/=Q^?g99gROe:ZB,[4,T
H+:[#:HA]_+)g[3V?&MV8W(,g.E#Nb)803.bB@Z<>V@/>91@e0T#9H7We+K6^84)
:8d&0:\8<V+NJ/-U<bYYP;1[IF)b17QEDC[#;Y(CaRZ8Qg+B<5->b,/C#b,L-F-_
/6C;XdCTS=UW80RTb+<f@(]CI_EF.fS/]C3a.9[\G<DD(FF-,PSR4Pa>U#E#P4Y,
ccQYA4f5Je?;=&X+_Ka<3S6>R2@ZY.T)Q2T04+b<6T-Y(ff=HIegaIEG#=JfKe^?
c0CG=OTN>O(ea2G^UeN47TQ4gV-Q?7/,E:>a,S1,>XacTKO2Ob5,c.;fHE0]N66d
>(QC1MY;]f\^^@-UdJX0[603KJBe,d9VY;Y/?A/EVWe\.]B5SWD=#F.aBOE[\_+)
;/E;RI]/T@@_2.RRAO+@(72FTIO--<104YQ<SM@58S[IHgJGB0A#EYWdDbebZR)F
\#>4c+^\JBV,RV0N+Z_>[O-(IKQD9[>d4X4)JGO;0,e[.)RJ0HLa22+>aN.N6-aQ
X>:-c0)26]8Zb<VET07LKcO1A558T-\\<F/5EBO)?-I>=L8;PcS6S=faZK1)1HHe
]G9AM5D9N_=b]38Z^PCV@1DE0@,@Z:I4R>Y4YdCI;A?>X..E/Z-N9<2/U?#H6X56
9CV.K;F#IdDgYD6])BXF8(?f-W/\)L^-&B#CbK/.JI2K30>H/C]/TRVCeY-f2-N2
fZ9&XdMH:,PT._HFOf:D4f(:]1>6DTHBZM_Pe:Vg_,ZaY;aK6fB1-#FTdJNKBf3f
F67fL(B-42=C8C#UOdBbcdIJ4E=WT.HN;SL\d;&\EB0LRZgTQWNB114-HG?Z#W=<
28\GW]/-6&E_\/JCTC-f;>17)B/N]OTP^6ZbK=6G^;?-f:?9d^-8D.[P.=)@+b,4
9VB=#IEG>,JM]86fNaO)VU(GYXb;fN^;F&P8S:IPKNLg,8P&-)&MARPRBd27NPN?
R.[\[O)92#Fa_.^)93(>)_OE(:SfU#PMF(M:gO(H\PIeWS2MM/8c0/5X=+;&fcB4
aE^ZWg,[g#588TV#5&VbMN1LO1FbVG@YI3\/9Y;bW.[5-.ZDRP#2M&e=/eEAC?,[
K,63#)gbD13\fZN6TbRcN?KXEfc#XfSgA4L1c/T1&AA]Z708RLLH9:fG69_]IG2.
:BD4I?-(c2&.^I8^95S@HR^0@;8PXeC.9Rg_cU=1e09Z&A7D]HQ68e\c6Qe6W23#
</=3RQ;<ZV:gO-cB=+65eG_/df/03IfALd1JWLa+&+?1GIHUWJ8aRW2DD2;ecUX=
H;V46dBeEQU^SK162H(B5&X5AZOYIW/R2,>BQJ-Q)YLVXA9IS(;4@AKCVV8^EDRd
W7OP1\J<DecR\_8P9YWYMHdR+U?Ib/-aR#,7=M<X(WHO3+[&&2F0>O1;T5691c+2
e]IOgFMHD@/ODRM<Y6[[Y#:Q4-668VOW\Z_7b?<JZPdPJPfE.2A+]C/>Q4(Z)87c
B&1L#SF86LMBd6]cZO>KQ-=CX&-S5H]9^[<:EB/)gg^,+-)Nba:I-X1cOQaUV+-Z
NgPb.f@1df.FQLfGHV:_&6He/&2H8f\ef9K3U(\8JMF0b<1P+VEFG5;9A_^EOc,e
NPC&PBIN5SYcM<54&J@[CLUP:L?3MD7/G#U<0L>C<A1.D?\:P@?:1g<L;BHd_gU&
MS=\@<=GG5<BBN>_DG[(4UC#/>LKOa]GZdKdRH7/OF5R(#4CG62A]97PN8F-C:U/
CF?J<+-G(\UYg/:N=;^4^<4I5f#_+X\HKeB_R+A.K>&:4STNIf51\f70:AL/[^SW
Ab4,g1O^4_d-V1/;5EP\dRJ>>U+C#SA4.=^-QLZHA\?VY)]5GGG(g)]ZHY5[86[Y
G=EX0\\BWL@TE6]I0Df&A,&D9]^<S1-[OH24SN/6D,)RK6Q/A)D[0Q8DZg;C\@07
)/>fL:>PH\Jb77A1QNF3A4c>DM)>]&4=VE+K\b20:AD_,-5)ZQ?]1GL=dSZM9g>e
P0OHG@).5<5NJD#fF]+68U2.0e+I3GNLJ@DF0[C[Ag_5F5M8O?9ZZ?5;DgbPQ@dA
5,8Ud>>1LGQM8H7K>PG,fS#R.OH<L\I-Of/TKGTLcQNC8;?M/]GIcFQ/4g&?OP.d
FS,)#g^EVN&UKYC]eeEA>77[IGC\TM3T_D,?FIf+NF+<#V\5)\3.\R,_/?Q(#E>H
<>#MFH/ORMK@]gW,XO9?7D3(I0,4V)g?83Z@>U3XP<.MG-Z/63Mg<&73/WQAX\Zg
;d=VK;CfJ_998WG7LSDe[OGZeGLe3JccT755A+K?]@R=E]L^:ONATGdf]7J^+T)0
+5>PFaH:TIZT/+A8^gCI43ZCdXE<Ec5Je^-OJR::2M0d??Vd&?3aDY3P^FTc8BW<
^/V2^_[&WJ[D9X^MUP?1D#LcdE2_PX2&a(H8MFQT2N:W:>E,5H5X\Yaa:AX;d6)G
HF::GCDB/FSZ>=7T#/J\fa:PXX^O9JB1:H8;YTLI^N6-BI=-HL-SGDA6351SB3,e
@0LKMF+67/>&#FU@=:E?_T5+?MfAaQB_/;J^RAK&U0[Za=Q?@<^H39WSV7_#NM1L
AceWGb_HZJ/NTMV.69I-B])e9U:/+.aP_>e;H&:0W/]V3d0JS4<7@c&H_KIK1[C&
SUCT/2M6L0O?0YfV(@@DVYa95(IQLgZOE6WdMeTeU_EdIf@HI)S?-TTAfGOJ=afB
I7d\;9LWCg#eR81XV/1I@GE;EBZY6HF2a/2V4UE/N)QY[V[]4TXP,b/N22Q8#FeG
.f>Xf3U9D7^6P)._B^GD77(^^^ZT:]eG(3[PV4aR.X(@]a-05THe<W?Ac-bLX,\<
b#M5WJZOMOW9MJ<dZ7NAT7O&9Pa+JAWA/][#^AZ)aG?)U(cJ?GGQWZ9.Yc,<S,6_
--MG.;P/Tb3JZa#76A&5RTWLN0[b0Rdf-1:\M?e=I9F[/bFcJc-=WUc)FTQ\&eR=
J_G)V-N0d&W)ZAN8)U6(]_86[/TPFDDA7&ARZb1TM7/,6_D+gCSc:]cL]VTJfI<?
Ka\,FR;8397CGL\9FDYFHK0&=]G:f&/E&:b6G@.B:[ed@SY/f(]#AGY\P00P,\VP
W@/MJ]b&R:J]UJP-GFTUGC3aS&MW3H/?N@TD2#+W7bC(55H4=34[DI[?F.#0]DQM
OLT(J)HL@f(K_6@C#I;YYO6E,HLX7855<Ncfg92\F0/L]9S10PFSUg^@RL>>R+&-
?;I@g-<@N8;AVe6OE;<_FA-_<A7.;H\^[T/=T5aZMG&54&RWN:M+33]BFZ23O-<A
KNMN3\##^VHQ):]ZK2T+&0CC^)gVA_58+X@.A:ESXK528/KEIP#Ead-UMO97?6B/
N)7N5Y1N^\06?5/FQd(GWC3(@QZFQ;Qe1E,&8Oe1W5a8c?^E/4D<TKUK_ZGZV8_=
@&-C,F\HU\Z8:IG-?1e66V@K7U/1V/.8U(5YG2#c-,@0/5?/gP].CLc;_9?)VZed
;96>,RG@W\J&_:V;IFWMf^Kg,N5MU^W_?)@>Y/@cB\?g#Yaae]O.>G_C#4G:_ZF7
&[Y?_^Y6ga&Sd69>QFf4HSc44(ZSIb>8GVXBcBf/>3R1\c-<V[?@UAf)[;c6&+&a
D)TNg90L_W.DIFd@f;BUM;O;/f_XP.Q9QV(cSJ;16e?XVN@US.#ZWb[EKH:b3,6_
WMd@9E=dZZ5>O,0/38Uc34.X1D_;E^L(JQ7VB#E>adCdNP#OX0HJ0Uc_&#:OA\QJ
ag/Ra9CM6MaED,b_Ge_I0795T:Ve\94:;R,b0:8.@e#AAZ_a6KN)6NHSfHeAWA>B
N<]WUY+d3#J9I7PH(YLG1VgY@5:G5:[0F>:6+SU6QHPI]\=Y:UWM?\N.eK=HcMRe
Qg71F^0^IbGW88I+\bGb1G-^Ad#XOg[4GJa:7DI9_9(^4e:Xc:8.63NfCCG@)UG6
2C.T6eA\=gRg[AJ;-E=BE^+&13:FT[7c,^5:W0>D28NReJCSW\]GZ1#=_/6:G[&A
5/-O25;2W<)g^,H<Q/(ACC.-;FdE)N,:;HIfI)E?Z6JYZHV,W-:C&[T8X6>?3BXR
?]+Y_-,UD\\[.Bc2C5-L.G9.IK2TME/UM1\f,JfH)N7W9RVT8cF#?.181f:35KYQ
MSC?ECL_fcD,2#5H+]G=-I>:=,X25[3eV:1,g.9?RP36L6S>S^Lc^Y?KJXU:S@?1
425WKNdA]XdeK/;QSV.(OW4ZL\7<ALA;7M9:)\/<:UP\eA;f^e7L]^bX6QV>._R#
(P2MR8XG212_1[9c&9)e=4<XBdKE2?d[fH76)4QGCL>;XSP#AIP7+8aB\?KQ1_,@
<M2@2AJE39J?AUIOXT8KLeD99cIG&4OWGOO4R1eT3S68#<XB=;e]YNV#VH226Q[.
8gLeM,8()AD./J@C7MH@^Yfag)==YJM+&@K(&^Y(C)@ST[bSB5CT,@,#R=BZ3=cU
gUC70H/)C;\OJ3_e\&NALN=.4XZ0TTV@+a_-O-AB7J3R>_9->U@ZZ,FSH/Ja2WP4
]HZVKR1SdUL/L9,QbW/+2RU2G]eMR)AU^XfHLC;]7AEO[G]Id&G66Q#]:SJ+4b3)
=OI[8]RQ.6=6#Ye.Vf]@7/aP>^]=//_IN7eQf@2[NBbK(T.#KE4BR0TN/FcI8\Lf
)[BfN+K(\8;VVUPQ8:c)M?Z+Qa#4dFU(NZeD3G=aZMG9PDZ=^+AI])R6Z>[c:M8=
QRdEA^X3])+O[U#L76Uc]5N/MG#5,M;.[E#U[UTI,cZ42P]E#BCQIV7^OQS3F9dW
/62SMWP9+^]PL@QGb.LX36/S5Q(&A_Q1Ab(G_5;8I#=P)UP,3[V++O7@30#ZfSKX
BZ7<KG3K,Q4^+VIP:6+2P^GVAQ^BKKXMLUSTM?0<WC0G[VLZE-,aEe^]E>#+e_D0
RGCUfXRf\4Gef5[RGKCP#a=B&1TML.g2NB+4@YDV;4d/BCG:^8E?Q:(/[CX8aTB-
S17(f9_[M2:PLI<70YgN0O,+/J7[d(+20dQfCQ6I)^KWTHc8dg9U<U>;>02=2_J8
E9T7XVce@D2(@1>(;&4PB/T.U\H6+TBK@T6(T<75B\fO+E9<O?>5=@B5NCH6WFVT
45/Y#gGD)66.S8]PMe3^+/KBWOgda5KgKDWQ_2\)=8?CAS((7N1L&(dUWc8SW559
2-FMUQeBd0-)AK-\,-3QJE4#[\JaR0dR<=Y-9Z;K,PR]A844NAB;XLBSM,&HDbBG
T)NEFW6\FH]=2cBBSYHaT0OA&U,-Re\11,7BX)FbN3eK20agHDG4+V1VS&ZCH6;]
/2#O7PeRabb+\U2=6(2)d1ga26:.K>R:DH,+NL5:NB:B/VVU16b@K(S)G3RYLe,8
TJBdSO:b25:b6a\5.)HNe+WSMU[KfCdC^KVBY@K[CNQef<I5Q^)Ve9/_TG^+-g4;
CH\2U6(G4SdYGQ/bO]8_EAL1?0]@>]2Fe1?.DJZH(d+8J7d=932USH@NU,+/MZW8
5W/J3LVD:aKNgF9HKUPaHJLU&F5#A1\1d[2V8fMD<^F\QfNU@dSZP5Z\5-)SU?cA
>gW.Y9JK-OW+RBQ\gg,GA+T8?;PQBV>+=aUH?FKITZ;Qag3eAEgBX#^b(M78daW+
>#?<T>JMZSG0g_\1S^BM8ODb]F.Y8aF[:)D>cVg,H=g5P;48@,9@bUa+\5V(ZFM.
18,>MQ0SWJNdUAD9_ACBUG^T^QF\F<(9#Z/:X>V3#IaJJgGP:T^cUI[FbV\GNA][
W^NCBc<@)4-Q^2]W@DBPOUXN>G7&IQ^FGURMR:\XCW6JN.^YDYSQPO\)BVFZB-N[
7VUDf7?\5e6H;&MM.W(@6?:dC+1V^[<O45@8[PC(O5Z9DI\=M_/&ae)dDcO6?/\g
<&]^U[_TDe)+A7<<g/>:GYNcJ5gR/84IL+V\Sc-CgE25[dM,[@5]gTU#bJ8f4IHN
SF.d_4GREFb65O/=M]KKKQVd6agS)+a?BcTF-5+/4CK)4)YP_6bE7eF<dDUI40O#
g>^1;E\;be1\22a;89I5X(R1&^3C0OLF(3XLLg:G22IQ54NEILfI?QbGN2e=DF9K
Z\\b;=Z).@8a@f,@55[&2P;HOL:aZ^,^Z<L\c\LQ_I\DQ6RB)B+Z@C:880X>0M0@
)FdMUfDCN98,W3[6ESND?5cQWQ5Fg_W8L]N@,7M9H?+_e@@@,#>OV2LRP0_<fdL/
F&+f\8+FC\;>@g^C)/f)_U_<4RW/1&@ZKf^^=.C.J]bD][/93g6Ka.\cFc[VH[A_
AF,HD-SXa.N&^(5T0XS?O=06#=R+U6]f\8NX)09dKHPCG&^:#4B31)V9:8?aQ(HS
G9O4.)XMf\K>#>dOFI8#W\/JHdQZSdf?b)EePA::KE3&a+VD[+]fX0NQ@@G55WQ]
XT-L+(]]P.O+)_HL)18DMJ42^Ua-33FMX,#8UVX<(<^XbAG-PV8+Ig;\ZTSLgW=3
\PC><A79G:CQXE+b8@CP[K/^M&b8fTd5I5MQJS^GY+/WN_MBg<Y4B_bFTR>,_+-J
,;)5-Y\>ge,&g77UZ=Q(5+J>)7P0_gR>7\@U6;4-,8/B3[.L==:d1bBT&5O?I5ZW
7G(#;^7?aB.GD5K8ee6[:FeJeVS(a1dc0gONMa,/Y=8@Q[e@6XS8.L420_;0#E0:
c=L>)fV0_CH)FP0=EQ^KP&>H^KN9BcZG3eB7Zd@[c-Ae]\\&ABZ\cIgX3<.XYdg(
T_D3+?T)(C0W.@CG4d+]2^]L?B32&-Id_#T-64_P&6\D-FBA]CEIS0S\,IY&Z4J1
7>J]=&(1e46.UCJ1S?J)K;DH]91Q&6F-F\N9=WI_C=Gc;cN:bNDTS8HW7&O=2?-F
)AJHEN&N.fAA?(UB3+VZc7K3.M.EcSIdN_dX5:CWDfGWO(#C7)Fa833A[RAD;O24
>?1e]NKbG:&BbSHMWZ300;C9&X[-f+)RZRgKaE5>+.9:VT9+B)X1cT:.+9@VbS+R
e5JWd2/D(;C>;>cS341U5ORG(\DCM.V4@f)-X8O;H=Ge;\WT5Ve>fI1+9:c5(7T?
Y;(&4R(6O3NXBM1_+_bJ@OXSL0K1#;+#??E(^.B/b^]bE-3T.R^ZTdUC:YggM.)g
67eT.a_#E\gYY<RIPB6(PD<II(\b\G^#A\fQc)Y0fW@_7Y^&C]aDg4_O.,&f8Y:/
CcgYBC=U^7fB:629g&F;:\N.P,?ZH7IT]1)B16N6f>.K2DCQA[?VVPeQOZ27Gd+X
)-UcT85O<Q5:V3#8d?M3@3MDC0NdV#^UG+F;Z#\P-^1KbbZ)]#9:^UdcWc?(^0-7
ANYcX7WA1Kb\]850a\6Cc>N1;HA,)Q1E;1[RGITXG?g]9^c<f(1MRcdgYBAJC&,=
10/#<@2MO?A(08NbH\,ggCE59&9A[=FdWeZ@TJa5=.0F@DB5.^Vb9+BW161;NSXD
,..-:@[c4;,H&@Z86EbU\RBV25SKXX(0^5JELVa^_>KY)>C30Y)+<509C#gg\@3W
<gS]fPKS1bd>[.-A_7(D;LgMc:I=LbF?f@_;#0_5)QfWJH=C4.Nb52(5_bB6-:<5
(M?)0(R<13XLDD0:51@_B,T_FR7-S=38YQW1.eJa/RU#3-PKE^eb-R(4/B<2:XA+
b+K)^c,U1JQ[=U/\1WgANTKW-_KDFL9gDBgKYZA(1QSS_&L.3V^,e=d^D/8&D?>F
QJ;AGdaP=)LGe?Da3VMN_?#8<Ga,:PT2>Q+-A:CCQT6[PTaGG2PLCBF,OP[gZIC&
U\Y_[/]5^R\KOL:+G,5A2TG?XJX#?/2Z5]]2R->P)2Q9W+?24b[-GI-c?C9EeSN=
JZH9K>B<VfegU+(NVMV^(<W+GIaXR;=B5B+2]S>9P^+,)^AJbbK,aY1f^HfL&I\=
<50K+)?OOM4>4;:&#=N@LMSV/?eN1#/b>C/:[XGT>B)J]C[\YESIDe;K>6&^Y8Nc
\HL)>F4e5=O9-.,7E4[L.VOW];W3P9^>N,\=KZRb]S)^H3>eb#T\OU#cW::J._09
KdE()HNcAc5;d(2XE9dgDdc+5F#_L>f/B?cGDGb2L3>,\fT-XH>@GIaP9/FMREGV
R6P9[VE+>0+ROL#[<-HcHMOU)@(A_V_HS#WbB-[6d7Y+9UPVJGC&[N-)\?fKK8S^
fX+gf5>,K/GddA8U2D8abX3-2L6@U1gN#cG7J.5NTQ5c#:WXVbEGa[U4DQ9[/f,F
-(4<b#X/;MX7G\YdC4T2^7E<0>OKHYO@F#c3.Yg)DZ3T)bLMY(WL-I(4RdKU1QM,
Ng)\e<4129&0ZDNX>USH(Y8@/CEf4;R0W3bCE:/I^(.[:S2S@#^X8.E##H-eGPY;
.IZB_F;3IPKee^ceL4KM;A/6&RBBGS@_\V07N7>D?C_K6Z-G,1V-RYO#ZaU:[_Y9
?SaA]IaH:J]ARa4#QgJ0d1OMPAONX7&D37RWbdX2Q[OX:DL<?P,1C/Q/Q:_DTJT1
NQ&PYcfERIN?MJ:RUK;+Z3BQ..?bV7SNU>.e#]GFML2dF8A\P52:C=<gYY(Jb2_R
M,NN.\F=33.U5XPM.R/44^AN[=a>_g?V-fWD?D:UfO\aXM>J[C;Se>\FN^1307^O
gA2Ce:/3b@g,U?X3\]E.O=G)E<5T,A,QPYDA2=G,4N3+NSdVf9Xf69&fN-7@Zf<:
/XAOdX;M[YZ5_2S<+.ZFW<.NJg^FL+__\V24Z.g=bE8(c6;F.#1YLDCDM)S,RS[D
<-NA&>T04<aD>9=dUX+e\28MCST4@e<>[^dRLUN)\=L_/PJGX6LgRHaDaf9b.S>5
&R)/Y=>:c/L.KSJ@?W[B[/CURcJ_03<W>#4c7#aWA\c=F#:1B[d/[9Xc^2/dV;1.
G&-13.&@a7(ebC^I-^0OO;28M_,83e/6#9fVf1DUZP-d)JW?]UBP8K[gfXBN[Z,Q
cFa,Z;Y=)E<@=^U2S?V;.4&#NDBYJZb/3/+?@1T>A(;7XZeMb@Md./fE^?+_E7]F
=PR:?:;-(Qbe-/b8O:fCC#78#GeJRJMgGd-13ZXPYd/H>BA82c6dOYU\.(YQ,bdG
La2#<4<N-K)gb0Se_7GY2KV&R-O;+T262)^QY;O,0Z5X.OD-If0>+.XCW5P]Nga8
Z9<CG0U+S80]P^cA.AGF8>7@S3NK71X>C1(^\:7+dK9G3,9(8EHc=7[P&E,^.cB-
\Ad?&_QTfLCV0.aE[#gOU/NWN+)\6<IRPXQD2\JNN8:#eUe[CY;+B0?[H-H?OD:#
VTD[f7.WG<PMM<2AGZUWCaDQ#2R5I:R2#CZ#]ZM4Y<Ba;S@8ZDd<-4H9FS\)cM+)
IDH@S6:)L+:bF/3TaeAF?>XXSb.31USO4H]G;+\.U4\H2QA^gQMf5()(G9H=VE+7
XVESBe2>+[2J=9>4XD^RGW8]ZOgE\WJ:W:)WU&9?J>c?(JC_dFI.]C.5>+HX&8BZ
2VBWH?_?X/.dEX-DPOW#a;_EgL2T=);I5gfbHRJ\/LbCVecD]L.U97[06Y:/&YUR
,g)I=:C\A#R-)^XPE:_F1[2Z8VcCfXG<IedZZ?:Z,C,<K\bQN2IK<^H\715+ZF\G
RM<gWRE/Qf7-1Ag4IEK4AN1O<f=(Df3;X&VaEd8OJUK4Ub>(]FK\dM?)B=gP@B0)
WbU.)L;WX]R+XIE_GEXZS50KY;a&D_3>[g4TBb^KR(Be-<OWf&H)QS=<WA>C58FL
7a-YII5[#(/a+)GeaO8DOT:8Y/Q[K=\H:06D:5SX2XD3;K,W=I,B;Q/;.P[df)BE
3_Xg__6,&6#[?d@)4bW<L1/VI(5:[?:A3TE]T=.4DL\==9-S\7\M5[3(IU038FPa
FF9Oe#4/8<2ScW4<E.;:Q^EUT>/Y38J\\U^+e[@[1b(Y@X(-.EJSCJ8bgDAXW;EU
GEBF:dQW>OGZ_(@0B/+Q5-Oe&V2/HHVVg1T1#bKC[WI91\(&M+<(K:J,5>9JM+>>
X7@IB&]f6Y@A,4GZS[#2Z&<<bc;e0?1M=-OX0J@5+=N>a.M.\.0);56GAX5CcI(R
F4IHHd2^RN[/eRcYTQJ()<+BBff>Z9a#+(IDM6[0JAeSI^AJ3gR&RcA2(D/^U^X<
ADgALW1U=+_.Zc3PK[5f?;>;2?-_5Z.:[@W6\)@^dKHCeT#&7^)DX^_/J[]1<0Wf
8:TDb,YL^<EQL-X7L.G9^?fgHXNO#EK>+eY9E&VDZaEf61VDg-NXL+49TZ&@5T-3
Ae^JLWA[KV6,Xb<BWDaag?J@cPX.fYc>U[2_PXABYce]XN1V//;(_g1QLEJ0L^A1
PL0Ad4M70eQgA0e)a5?#)NHG(Q=cVe?1M\&/</6QG\X@&:YWK7ffH:UgWFP+9,#Z
^;]=BPa)I+Cg)9R&6W,gPX21)=(&D(34<AD]E9_(72KU5J_)@ZBEcI5Q@\<D_4ZZ
#V6CU<IcUbCBYa<=&#WWRGg:1&MYP<fJa(a>(SLgJA+QQM@:<7Y:=aWD#.DcF1MJ
[bYc>CG1D\UHAFS.=C;[NB):Ie;N=F?-U8H-9N8WeU[+4M5.B6QJ0-T6./+M(d]9
#2DgIX,8&geH)Y_BFD_+YFA--9;+R:8HY:^_HZ]E78QS_(Me_>(g1Bcg6(^PPUKa
Be6=F/6ab?PM>P7e=F=&;MXEb)E41,0Q8+E9[/aKVb>.?NF[H+>dfRc=[-O^V3G9
X5^H0JDP-g87Y5?DT)^J-(HE?IXP#XYH<=SXf.,BSZUOeEJVQJ/fOG1BN0#,1/\<
J^07d06DFVaJXD[FSJ\<K&#W#3>W#;^QF>_X5V:.95[T?.M-d#QIL4-O+:5N+S]:
CL9^BJYILQ2-_Z0M89ee=Q8dT@^H>fF/_IW,@5]5DbdBDXf+9,G)3C_0g5e0/^YP
[+_ST#]XRdKTY)QD=[4:849d[,7\)d&PDg^F5Te(HDgD/VC,H)5AV+@F;g/&6QZ[
cBBO#3+HP==)/YO39,#.-M27)>9+/;I4Pc0QaI<fH3ZCUX0bQ\9P)5a10g&W1)Z0
=KQ9H;?]dI>]VT-WaV4b?]eL.;ELT(#:FS163)@K/;JRgKD5PIED;\HAD+98FHd#
5S(Z>3TU^Xf)I1CA=e-5J]OdIQ77\5g96Q3__/8065BBJB>EIdR_9RR.ZIHCWf+9
@-b[aM\F54RfO_F9N>Q6]JT><N(@PIQ6VJFV?:5WeQbd)8gK0I2?)Q-c5#9GJYXT
I=H)C==XEegQfd+[XdYG1(XJZRfe\Z)DV;;QKH08cGag5-,V.We3U5)@.ATOJ(T7
V[aNZ@AZWXZEY_ALa7g603+/6c8bW]gLFUV_CeL#FEWf\RW.#:g2782)(UL8PZW?
Rd@R]T/18+[_RgeX7^-H8G&P<b6A1V?F]cfXVI3#)/K:875:>GAPU#-Y)>10N0CV
V#K@3g=e/QXbIK+e5/X#XM&T?O_XMH^/[:XJJQW+f#0[XGVRED8Z=)2U0^D7L8/^
OS4ZHZF47>\SDN8ad_B&7TY>\;:?(d(CX&]K[20&^6KSaR)f\If;,&96W74]-8TD
#DRPJF=3[&=Te6;C&^0AWCgJ&.7PWCPDJ\QD/85(60SD6g<caM95-78DF-dF^L#5
L4E>C7G\O7f2MKSP5<UR>_dQ6)^V:4U>972SKG0QCY+d=8M,BZ@J;RT:WS?.E:5?
d9S:P5/f^fA6.g&)@/4ON3Sf<JLVTON1L#X=\bQSG&:3EeXKf)6LV@cF(HVG=\f<
MZb<6N^Je.Q68&B6Y])9):1]085Ngfg)]@_B:)07P1[;TBJd8#HYN7C?RWaAKSdK
Pa?>DVe:F^717P_41dS)(JPZX76?-Q[eH0d_6R_?b@-5D3EE\1/?\?X)SZJ9FCVR
a5:E,;:+eOY+(bYLBR;L?5(:f+&4H\WD)\R[^S,W)=YKF#-50T]cW<,6VD5,[7d/
R8]K_WaPBUeF\CBfV+;1QTH70HI#LbY4>DJ/S?V:aMDE2e2VDe1N<.bB?\^1]dWd
0GX1Y9c<VC);>T<X<H2?0gEOH_\>6^QcREIHL4dA^Q/1W35?NgH#](\f?D\e1X<=
-B\I?AB]]UNAX^4^5_=.92aG:0gb?5-\71367_42YI<M4;=e]gF+aTeX+A3,0O[:
)\[(1[P8ALW6L:9&UKfJ6Ga8SOVbZ:EaT8&_b0SHSVK\-U83FgTL)LG+eBF(V8EX
\>?CK<g4Z7d+_2@IEM3)fQdP\R1F_2:;MPZaHG:KWUQ-Z6>,J1R6;eX.R+_1[M08
Y+Ka@[B&<N+(-],eEafYACV]+_^]W/R;ZWNOdSS^[XVX.[GeK82@6_GZL>f1]+HD
dBR?FMU_FGJccb74dRNJ4UL@:AaCF2&-ANO3gRZDV4EJ@c-aV:82DJ;d>.YYP(EQ
[RJ_(8[H5e<Zf?fSe/6O8VSZ&SA2IA/Y+;+:]?gc>9RSEBSF8[1Ab=HTH4XRLI9G
c.I=Q#MZP+aX(C7S;34&58Ff+PCNfR&9E0H6\L<X[e-[C9COHE=AW5ggQ[(fgD)O
M<VQP-IPC6A-L=Md,KDcE9PB<O1aGeU;+\I-:+59gNTV.L21KCb&\dOC/>SYD/bQ
dSaH#=g7\CO=^2\F=37:^_+Ne>GR.1YZ+Hfa[7ZNaKK8RZUFXH)9+.PB6<C_(M3-
5#BPE2_VP7&1F[OeYWK\;gP306@J(:S<A@#ASELZF6L[L<MgAA3CcX6+S.CZWF.I
=8L<;b&>Gb)0O@FS@#XSW1)W-BF3<@+&ObG#\Nd[NRJDUUT]YNPge(fOM?AaI\@K
1SfV.BbAHY=JNeVS@g?YZbR6/2f@?Q#b@BaQ#-Q43Z/&2Q(UUXY.I/(=M\U,#FdD
9(HIcF=>?e_MQ9HXO7baWd536L=M]1/-8GVYAc\6eS@3b(8Of[VP2eGPZ3F=D)>-
K;B+NOB?8J./;A,OFf5VRA1):PLUK=?IOfOefW56/:@:.L,F(\@,DR:-aG019.@.
5I-?<T-IGSZ2[03A4J\)ATM568_A19S,UE=gT-F_87ZCgHL7a1&AD=a++g,#Y].P
[):ROK--20]).gg[=_fT,>FM1e[fR[g\3(]9<(22gG0);_86EB=;\1HeW>g+TWa=
X4<d/\^)JeSI:12N)eMH8)-?PL(F1:1U8IHTTW:e([?b;aAd?)4\LC1g[]B_VMD>
XLg3@Y/FV6<D63#&E@9.[7K)1HLbS[?AdO?8@\5=^Db=Na6?EI0.0b5fQO+F\7YW
<cS2(=bZ>[;.T3TeWW&BAX1/P&/>?PM./Y1F-W83)(H9SXC7-2KTHP=\H)#<7MaS
_L(1_F2NUe@K^d>_,Ld>YOY8D=E1);@_B^H&M8ND?&G0@.d4S:G82g5VZ6IWdRI]
]fcMWcY842&QFZd0@He08\QZ9XRTS(D5F=\//ZB&0FCC7MU?W=/&3](ZGLgW[VTR
.2[0,(Yc0)QJ[d2.L5F=1]/8=];;bXZ=Hac:J]&L1;S0c7#T_dYBa;N\PEVQ07\V
NC;EOO<]PJ@eBe^2VYJX:.]IXG\V\B[=OZ;+KW_^X1-f@TX??RWALfcPX24SI]=I
edH6H(d,7EVMDJ:a3ST>:)<>>d[)c7T\Ma^B=ee8@F:)X;:F;)B3:#3K5)CfVe9+
fNY5/T7J3E&]SGC[6K0Y(W@N@1N.LY^30)/ePNW3@+gQgPE^J-gP(C3J[J7QH;WU
PO>.7LB/DB3Q]M@2.D?Z.LdZR;(Xc,<KH3f]fcU:LbQ^91]Ib]>\[8[U\Xe0[_WP
X<8A83a\K=dM>EA[E@]\0:B:5Q^42RBVSBP]VY2UTF4[Qc];+Y-E.^KC-_a_8)B5
eHM_]6U\^;Be11a&,A.H3@A#M>ZJ_1L))cA&RKL?,7(9Lded&F@8g4MT65^UXIe,
HM<IbgF]?;FBI21)J4,.YZA)XTf7g.;GVJRXd,>6,Q6OT.IQWB(-Mc_<=B0aGc<G
cg<G(M#ZgNODfF^IJS4&_1bHH,GS69A1./\P_SS2=cKCZ1[^^Ag1^Ec<9&gLM<<7
R]:(=LeQU@F25^C6R57BFDKWXU<b@0TKcf1c>5g\##Q\8]b3I1,D\/S51_&6JQdb
[Z1UU,V&=)af=:[0HCI(4(5(b;UOM?ZB^JI2f<YHBd:8M2RDZ->I[.eSN)QWRFed
I:67@5;-MMR@+W_6Q?2HK,c]=,/aT6:cXRK0MSgWc&<0N51/<GSB_V5DA/aaKU,Y
L8f-I@42Nc_.IDE2\Lg+PFR1;V/+5RJ3N93EZE:]Bd@A:=R\Z-C:959>Y39<FM/I
/]0gc<[,&;5=(??#1-V;K[M2&b95X_==[ca)3/,4d.4Zg#(8#&<a^MOb3G&>fbDD
Ia4eZIL5_#C]9G08d5Ye>S[8\<cYbIaO7;_6G(KC[@89W+AFZ?+,8.EFaT[TR<IL
B4]\-Z/+gT64(-A0W&V-CAf23I_ee,D-EH61fLKHAgG]DGMKX9S)L-RF.]gLA#8-
QfQ&;VfD<S]de6J[B6PHJ-4OG,\7X<0AJ296N5_GA]O@O[VeW/HM,F>@HZRV];CM
8Jc6/Y[GZUbIBQTR9DB@1Xf20U?S0L)A&4LQ)ANRO/=W).dVb5)8g=?R?;HYbC&G
Y<K#1LL57[<LW-+M&ZfEYe+F>R:,]TffM59@=8G?PO@1()0MEAY1/3\+S7.1;>eB
]B0<+OK41TaO(cZdXe@H@LFJMe/fagGeEJfIFB(BU8ea&bL+IdUfFL]Q+b7e2Q^J
M)=JJZ>KGF8X;&WYM67:_TGeIeRVfZ;bfMW+.)/#H;^=ab3WL,ge>R_1RcWZUG)9
<Mc3JBg8?1Hb<9SRPNN3Z#<]KQ2@/(?;\&5XZF04)/.#DHf31;Q<(I<7V6;970_>
X/H[U4?X+Wg^2UTUS&<2ePW:;K:D;^d@MN9?;&?2SD-YTee.LW9&X(<\8+8I/TDL
KJ-+VP2D0@21>ZJA=UR1(c.?Oc7XeRA</Gc4X5:DD;3VX\NH:S^(1K=[?-PaUgM@
+CCOQPMf]).EfU6AeKgg8(gD8YX#f_J]@4[c^N+,0<+dFZG,TW>cg8GPe3:.@RXZ
HOIeAc^Dd@UT-aI6?8aMAIEZ72S?9Z(GH0^<8/:6\+Y,7/F=F,aU1ZR(@EWQbB2F
FfF#H^dVEM[>=L057@HTf0QMYN?e(]4G@2QGb\FUAN\4a>M/e.A;N5f97^7eE6[#
De>^-^6-eaN366.b4aX+^=G:^Cg7?U\gf?0S]^Y&.MZ(2AYL:U9431K;XZ=[_T).
1agI,4-Cb;2YNRJ/L6(f=Hb]6^:Kf=4,P,_=VOJR<49e/e..[093D<Nb6,;?cDdb
-V)Y6[0\7-&0C2Mb/:;6Ff2S.I3865XYJU3eINQ@B\A-e=V];46U]U,cDX:SLZ3=
W)J#b[;+8bK(Y+.1#1P+Vf#-X/TgW[,c5UBFeS528+;X<HIC05&RN\:-FaNT9;M1
gd/2fZW\02AG?7@?AXT=Be7SI]fSYR[6<;R?N](?[_Z4VaV=[92\f?F\=2,.>429
,F=1-G0R(24Y<:M169SBU6X-U^Wc0dYL-Dgc^Ia+X6)+N<5+c5XNM6Z:&P>D?IaK
>QD4[79)FI/UO0T78MfSQ>ZD+]>gW/9PeZ6bSWS:Q^RM+XL=1=c3fb52J?D)JKON
U?[^U/CUQ^P=?=C-4NdE-8C1(cEa:>6=XTL_AJ7P)14V-ZYGSUJOHLV;,:cQO0VA
TCBW38B),7DZcK5)3BCfUK+=?;=C>e3?0EHQgO(=>McA6X0MEUFaV<)J)&8/AONe
?VHSS=-,Sa=ReX)=Cf_ZG>IJg.I><9FOP?EL-0TR40#\BCdY^[T/,d^Y]OML=U=Y
.Pg,/OB;B#&&R52>+c;]0:^TcgQ^:.BC/gQ7-7A/\b?@W&c_c@0/)MC)IYP10ACf
Z>[(#c,P>&6GG<2)U;J0-I&;@5QE=?G-f]VZJL-4Y\5W/<WFHe[JD;9#Y\UbeJ2&
HL:+0H25#W8Q,E98:^5[(6[P(_J\,XRgJ@&VA013d&Y#P\AQDQEac0WIQ/A]22S2
+^\d29F5PA4c4OK8MT&-X,TIQDDe[;0/<UOQ_:3Y=PI0ST&_]E32+]#I@9BDUf&f
]eBR=[I0eA/R)F8B-PJf1aL^,5T;g#;HRdc0GU8U2Z=K:(ZDP\,0BHf^[B+3<[,W
GG>bFXOgX13Q(bBWdH7KF@<)WN=,dOc<BSN4R73FIfL>1\eD?@S1DWWNUY1EZ^UR
WSV\X[^C1H#51.P[-(?Y<fQ8O121eR_K]NB/>HTLMHV:YA^=3FYJGF-(aH/I/@OT
2+,f:Df0ZN_>d4[?,1d)]3PAG_<[0<^VC3>NN]aS<_9H-3c[5[H<DE2]^R(,g=W0
]<UB.^.;<MI@F:1MNg24BM&a3XSOLbK=65:#2/]@g<1<PNDVF62H[71<6A#g63&N
]f5\@dSYCXc51G(8BN/e1)9]2P,]1g;EFL-Ie6)C)579LNY&ZTYCac4WATd[b__T
K[1WH,#7+D=5Q1Ocfg-4[_0]+O5aSD)L28PWTAHg3f0fU&,=R+P)1R;Ya2W,F]T_
&^fP:I\J][<)22+K^7S9_,S]ZA_Y/fA4gNB)LA16bL>KV;3@IB9A_2U@,(1/[c\9
Vc@>=2/9^7)b\).;[[4fFMV8_2aL.NMN^d<(3JZ-e0]N=Q@Y/X3B8If\5CSZ3OHK
ae<55>GNTP.aLZYA(C/V[B0^)TZ,aU.21W8AJcAH7/LcS.YUWE5VD#C8+e^S9.>2
P?Nd;CY1LSJBK1e_;Y6H\8T7HQ6?@.8,[HVJ_0J:JJ+/[8WMeFgT_S&Ec0(Q05:d
[;VFR_:L^-K@J&=R_^?/5XKY)[;A=8PTJ+5:?D1QA-Q^8EKJ2M9,^CY4<NED14f#
:ZAI[_FL2)OL6:/]==5cU36<@eDBG+2Xe3Rc3[9e(A_#:)6/S5ONSW+)LT2Y/]#N
D&,9>cL4(7?Wf9GCa^I23gf)F<:4EC>U+ARS)@J];;GLcTKD1/YdY_[T?1@3BX+U
S7=R)/d92WTHDZFM=T89:Z&E5&:3YNK:\9)9PN&0@\@;5^<B\>^b.Mbc=e1]0H=g
e>SGU>S-a.?I.CBAUASdd8b&.8a6:0]I:82]U-5;C\)[]=?4>Kf0P(\fYW#SGae5
L_4J]E6^>d1W4&5F_P_dWNN8PXLU#0#RESZ/+^51-e\ba8fDa8M9\@U:JTdKe=AV
aC?Lg/=f+VFaZA-/?6Y9c:6?V0&Cb&d)UD@GNb)G+aVdIIFH7HRR.-_]DTd>2+#1
PKJ<QVR#D;f:8b9PS2(MS331M:Z?6:,KIAfPee4a,2YB_;0(B26P]Ye7@:1^1QS=
WOR0V7S@4_6C4&3>-.RW2JW3]I(?,eH5+CF:Z9_bOYa;Z>Q&DUJ#.d^Q9^S=[S]4
HNX6c2b4AO3FYA?=07Yd,WF#d=DG5&#_g4X^ZHH7Hg:71[1Q^K6bKBI_0@FQV5T6
0#EbM\bBJE@DKCU?U]623-L.eKLPCG:Z+@O-N8UJG(N2(:<M:0?=97.HR++7a1P4
[LT[(WX_gI[K8N9[bP+ZG,X<-;+REQG=F6@>WEIQU142;Da#HKGB56\<+WbMJ#0e
PZ(a+]C8Fa8QTS/:@B_QHB_#fYR\EOAEQ62:1]8L\c?/6L&SM.K@\#?FY68[G_&?
9_.f.;,TIYf>YKS[Yc+4JO4;:b6W:,/9aK111YT^>J,6MQ<9;f4PVIT,:\99_FI8
&-LU^@Q8\(._Z>OHW\fgTPCP[S,.-5Q6VT]X./[:f[dTJWJ4N08L<3cCD>6G0Q4-
0R,d7.Q),&EF6X.e8Wa08ZXD;1)P>F#:HNWb?0/1\]S(ab#HcQ:ed2Le)[Z8]-@_
J5PDbfgYI1J4<g0R.#bJY,(+Y&W4W0.J7XX6g(SU+74VbgVR0U-5/K\@<>U<@&(I
.<4XVEU/-R_U2UX6-L]6?QI?IR:3:2&GNc9<.&HUL)U8FC6JK>5?>ba(^.(?eX=6
6Y,MBS@gY6X28NYVBJ59;7ecW]cAK?8Z#TP2(46\bYCdPLO=LQ,Y\.&@H-bK7_bD
e.&8QC+-RU,;C,.K&^b8I,eBVMWOg]gLNC9Z>6)A7O_.fNA_Q+Id1F_&?HD=eD8H
9_Z@Gf0XE8NYY,eYT<7&/BT;1AIZ.O]9N9fUcL)G8S2D/RX:F@6XXL71L48Z3HUR
/Ha5fH>1?[;dI1EcP.3?:f&E@JH?DZg-)8[43+PJDTHZ+S,J^,-ADfMU@B+-0T=E
Tf6a2=&Y(FIXbK;-TJX4V0D(,=^AMPdLF&FHH:;]SSVP.d&72^[>];?agDcVRE\O
5]_(?a,#LfC&g_SGY.8>DbPZVQ&QdNC)023Q;2B4O7/AdC<[#\dGS/LO2fNa+g08
GeZPg8IR[THN(+)Y2a/@dV7U2;J,=2Y&,1Q#XSND5f.Tg5<(O]7WcLCf__MVN8]J
egYB?(0CbDc&VLE0#=/._^22TXF5=.W&L@;g?Z\[0#=W<Ud:S,L(eK8>T^LKZN+U
GKQ6AX;NA4SF<e3e=_L+L\?OL)\&/M7H-K_P\M(SFe<JR;B4F/ON=YacD_U]C)=)
&[GT:b1B?YF2<7-=\b03aTFX4W)gS-)/ZB>Y#1>fAS])Me[LDfB>aM3_R12L(L^L
K7W36(6bV1R1&_/<HS1?1P_bWEUQdb4&,X/,BG6(HQ[5GWV4TY70:=G72V=.)2K,
d=.<WdeYa>[.:):<@&L:J,,ULIe=+-a&a39HF0MG<P#@)8P8<CR[^TIAK-&=)Y9O
^785P=^#T8_9WW=:?<HIIE]O8_\4Lc4E7)PW;#?Bd]S79,1Bae?WeMMN>M:=[FL4
;bY7EYEa8D7:<O9,10NC//>\2,EJMb_,I/SB<Qa?B=#dR<?dD()A0G?Ied4-e_67
U\-MZe,(R#L\ScYcVSOVaOFDb.UE[,/JKU]FL73#CTI>g@b2DLB&Qf<X#FZ6B&U,
7gK2f9PRC(N2)<^_V,2MJ<K(([VFC4eM&SLY;Xb]LJ3FTCb_X2Q6Y9=B@\F^#I-\
4)8#XEU7H-Tg1Y/2W<aG1:LR._9=gP]<)(>Mc>I:gP51:=7SZKDQ(MP/X;5dC162
^8446SU^UO9H(S.-e(:\E@c.gN=_R7BD1AN]c;gM<^O/:47[eCBXKE)Z=9B=?]9^
YCY6Q=2-&?;JJX/;KY,K@e0JH5>6D;+PS<BDV[OH(,L_8<8,0Gc2E(dYCcCA;0JX
0,@V7IV2==WGcEO64R3P=.<Lgba[.JQe&QNXG69UFFfC\LUe@),7(0+=UA,Z\b[A
e9M:#b6I(J+H9f@AK0,NdgHbgY<+Q=OWJJVCC57-<G2AI&J?JE+cXgY_419_J,^/
^Q/@GU8R37DUdX.Y0;7,\/-Oa7F,_,E<D(>QYX3ac^e#X7^VNLO?>FX;Ub86KJ\f
a]dKY3:+C[OI>I\=a0L]14Qe4,-9IMSQL8#3fO^_F?A<RWA0R2:VV,XP;\12=dXD
_>[JSP@4(6H[[4Tc0C#bW#R6TIe?e,gU=Se,U_X+6Iea0L<4]-D7;6UMc;:1[B<Y
4/;PB>-&TV/4fO@MI0/.E4JQC/4FO=--:N0TY[_/e8+g#cO1-\,-T,>BDVMg,S5X
B2:TT_/K?6?dM<9I?NHM=d]Y<bTY[1fU9MQ4>UaWX]O(PN7E\g[CG;T^]UXZ:\73
@A8DcBABZ=UR<ZYg=DF510d)<.XI/Z)I;+]TC56@CcIZ:[d&bSAG&Kg&S\e^?a#&
a<PEb16H,N1LL7@A>4A3RBTaLUD@6HFUK5AMMWT8.D<RS6fEBcXAHaY4)OI\2B6D
0ZNPIg(@f&dK:_L7U-9#c3(R]Ta^8)>O1Nd4X<U:/85#C+@g9gQ)G\]73O>5Y1UL
bTWJ7_5gB:9VCWCIf/)G520d(EU[.4.YgES\@3=UdZ1U1(4_B]#-H(gBba;JH\:_
KQ)V?EWE/JT>?.\ga;fXH.XUA2YL/]dW1XR5;RLS&71R3@g@Z>I,=(>6a&U.VL+?
P8=WK9c14PO>eI##e0^1K\]&-\W)7TOce:fM/P]K?,B;)292Pf^/-DJQ1^O0U)1L
H3DfGBAIJ?dSbL6c_35X3]291IdBT42OL[[=9I+KDeL2)/XX+CPbU^2<R7e[FZ4G
KA>;Jb7a2OX/(?V.N?fAF+4-XcDI.E^)VMLV+YeJ=EHgb2G8D4)+cYM0ST@8F6+8
JO=@cJO:#H<@HTHI\6OV4Zg6#E/RUeeO=HXXM2.gY,<c7D@Q_,9@F4KN?BN?I=>D
=3)@@](<?[;,=gL1EAN(DRg2bfOU^GXABbe,[E(UFN5=-b^f-f;=fIH=(+@fB^c]
1<&eg:LZ<<aG9EMb>EHDNI3VU:K).WLW,cAMf+D:?MF0e;]0MZOK53PR>?G/(Yb8
W&\=#BJa]\QW971:&&Q?)(UCHP.WB=EM<2-+GHeK,cXc_[4,aV>V6V^/#P?dV/Y[
11Q?G8eKL=A(4?W\U;@cV5=:+@9<3\T-X,>FV&f6d_W^^5aN4S0L8^-SG.)M2G[Q
eBaMVeSU+I<2++Wda>Z=@DYg0)A2S9CgB=1?aadaIFIDcH0fZ4N_3K9(G:=0<^d,
S:TX6-/>\0<e:;)1aQS+F:eV_aLK@f2MJ.BMAE-#&<+Ke[A>S;PLP&@,3g+J5H-d
0>g2+:2)S7ZTSF#[dbTgZBBHH(Wa+.7W9gefZZ\J0=;/#bebcV2T5O_ET6=Kc3Ve
f]UEe@1CKcNGV^2?2e#Md,I1NYX#4cY27\YAOPGB6)5.?J?Q?f]6gGA)&=.DP0T?
]7QS#1PS]Y5KY^4;<7Z5V549-&R.c5+eJEX4MY\V4AA2P+2Eg-EE?M3B2ZZC4NgI
_DaGQU_RD)C3<^/H\UT\.<GKcY:E^>ed82H-VL9M1-b167+BDFdDGTE-_275&VZ/
2/].:3V&3;>J]+Og1C9^)Z+.6SddJXOg.<fd.+QNX7\T[)SK.:;TL5NKdA.PZWf5
(I_PU4?[DBdZ,HTI.;:E<Ye-YeM-WcO:(Q<8Q/aHXgPd38?aZ7G<2FMGPQ/R6XFa
f?ZbFOYL1CSC\M4f.a\aNAcJLUdc2+a/B/#B.bA]E]8Q3&1g5V[(?GIY<fLWKN79
g-/(/#[P021SJ.YeM4=?cg71Y/#60VGXQgf(S8eT)5A2THZJ1Sc@19RSKAD]g4c3
X=Y=[PM\(E?9c5fcWXgZ#(Q_cg1HNJD3<T?XQV0-\LNLU)g3Re/1:10W>]\87_9C
<7?g#2U<15Q@5EbZePbQK6V2+O4X-XN.IHgIPR6E9d7(]W^VRAcMD5;ZZ,J6-URP
]7e+e0.(cH?P9A4X)5A1=4&IW58&(.#Ob&gW_\XTRd>+fMH>?G>1I.TW86#1BW1W
6@I:?U\6gBQ:d.X+;I,c+cKXJNUOG]SXdHW.ZT[629B12[0[SHc[g@^C,<M,5TcV
7.EP2Ya7IW7d:8f0@DBd^OQ)VD90L^>NJ)fXD+G1@J/0&2Sa;-\C;\XaX?)H5TMK
&5BSSPL2:[J2gIdB^D?BL]R=7K(1YL<I+#[-W@A^].L/]/1XVX,_HW[KV7N0Z.1U
.?\:QG-(eO^1JHLf6GdQE.EJ)2KK^31R(/<RKKZCXf&bBP.X#(.41Xb7W0dSV)[T
5L3DfRMB^42DSLKfEa;RQ]MM3N6,;.<JL096cI>g.ZQbdbJ.ADIJ^f3=/=[2L6?g
<9\)2Y]RKD:=bU0,bKQ^<a+,-QUP)0[a,U)Y14SId2[M@[M>TD50fZ1KTd,_E.N2
+/IW^KG#e4(WLg=+^]Va<2961/6DU(]K9B_2_D/<)(7c^UR:@LK2Z+LE^)];a;8F
)eA:ELdVeRf&2&^26X<6,C?F/eC3/&A1]f3,=00B=R;M0Z:+a4DPT/bPR=27.7K8
SWJ=_,)&/1R6J,9H81&=<aC+WQ@dAAJcR/Id);=90T.)F9JL7VH4-4UZDAPg9S>Q
&3@4O3)::M>63QOAgbGWMJ3=e>Z-[/eB<MLR,HaT4IPHZ2-OGS:&M;[(-(VMGc.?
2FS8#7R.:K.EcOIc_PT43L\W>M[b)2F5ZOS;8f==1MaWNXe:O07BKX._;QO5?YN+
G)>M9=Wc8ZD<.1<bcWJVe^3?2+e62AI_+WdCH?1J5LS&P9B\c:]OMVMfae\I=O1a
=,R46-1X)Y9\Q2E)P-C>;4U@-c>(/fVXCICM#N>6+<g(G7X_W7(0/F-[E>EY4^MC
Z0cCOe5SgZd;19@0d&4\LWT8G12/18>@#@\427G1cTPXEd<^OW<QL76d[#Q1K<S)
?P.<45FOePcbFYN85_QFDeI]C=f^SF8fVW-2e67R5MRCdSg9_^fK?]#TCb#E#2]]
_^eO_W8a,?P<D,I0afKg-cf-5TQ[4/W-J(G\5RD5aBP[KA,;Z&?L;MX41DK#G^<K
#1aB[Ne9cMA#:/1aUZ)J243;5H7/4^RU=]<;/[V)=)&DI_E@SPBCCFS-#68:8T]R
dRTdD91fdBFJ[+[TGO.K43UQ1_,E46KMe00Tc7+LWIXCd]J9,6YM_3\eAd)P3<Q<
48][&(+BG0.UT?56B/LE9f8fKU\@UR/NG@@f6J.e&AY_M[_FC[JXgFETC+U^M6dA
bH4S8YJ:1;g8#a>H(-8-&Y;<,R]LH6>49=P=OHRNF>@^&d\ReVd,&]g)ZP-^NEWb
9A_A#ZU2PJ?7<-+AR0)MU;-&YgU#T2#.#CD(RW<a>1I7AHSEN4KI8[WOC.J;76MR
;Oa4^8Z]G+T6#8(T)Wc>\XR8W&JH7C[ZP1O?GKdKFO[Ng73,^9MC1/VP)I98a_=D
4G.+#R2f0_KQ=JR12A4MM8VYE(.fOc-[,D;25#E327&LI3(K05SOU/<,0?8D;b?B
^;>f9TaI#D2@UUQ@=N]dVA8;T41f(c<[1E>B#TRP/H@&JS[]^G1S,/?QO-DcSK;U
F&C_/#AG<EU0UK)ZeEN8XP8A6(._>P#9HRY0#RMPVZX=M)ZYASTA_ROB=fObVF5b
5Z(EZX&gM07#2OaX5Q-KR&>8T9W?[fbPdKNc?H)2,M?La&e8+f&Idc)TDP)>b+#G
RgY8[+7f=EDFd]R?(\4(aa3<H..60?ZaU<:^FbQbc5=b1]7L54?(GZ.3OfNH6)PV
d/A7MgX25(g-:Xg&R?e=OY6QLTW\JaVZWLJV&gD7TZd)4,7<.^RW/d7O:E#.S^CN
^AXb:FEP;K2MXf73)T46[YN2&4S.0<Y[IF4Q:00X#gdR0+Y26d+\:>Z^14<LT-<_
;[CUR_C7(/BOefdJ_>O2:\O5P[ScFGBH[)@c9N#47)dCg+V..M+\f;@16YFg@.19
e8A&^M8+XNYf/Na^TMIKTD.<W9L6<C1KdN/?R(@2gfH=F..B;:19L]Pd9]T5cKDG
CY0>O?_WNMJbJT:^H.QBF.ag4Bb@]\G2)V7Cd9)gNSIR#M#C12aJSD&B/U?Y9T:[
I&MRM]N0/c]faE,3FI&7K1<9@g>UTQc]0^M10-97SYW,b;S8)JJ=B.H?<E&[76.E
@HL,_)&+/.5d0TgDNY/<F7JHE#WZ=YSF6(^C7R.;WH:Db3H0;;=:cBG/9OJ,T.cF
dQ(c&3Nc,J-M_[>^>7>OdYQ<1>CE.FT7B?Ka@1V&QN&Re7U+.B>dgT7M\1DR(E)f
R@N>a/F,7:eWb2(UI&A/IE3XT1-=+^R(Rb[Pf&7-E9ABe25K=AcX1T5GM#&b>4Jd
D807ICeTXfJ8a_64+b<P.Y0-K:4dIX1^gJe]1J4ANLG57J/36#=4S;W(0TbR(R89
88IMQX/K+]J_U2.Y]g#]P;ET[IdC7A4L@AUSY-J-\7^QH1&STZK^<?W]_4Y+T1TL
3.HA<gAgS_4SabA(c_ECeSa->FfT#W:&5N4@.&_L;._QEG\AMGBBZaQ3)(M-,0^T
M2DP&GYE#L\_<=GOV:C+HfJ,9)<>VXXQ_1LRN#e@-I-#5>WA#.5Z7,bE6]P<T&3D
GM\&?^2UOAN:^T-&T?BKM1Je4AddQEQS#0?XJ5:QG\?;+9FBKA?1X(HAWM=?S0E@
J9E./#;OJD+Ya>BZ=:cL-W2D:7NQ9M1,a3bSMA@6&WUY3L?JWQ2+#&RbV;,]:FB6
N^U34e1IWS<aU@Yf-.Ja-A/]>]IM\NXJdU);I(28WC1KVWb5\eJ1&(VcUPceN:g-
Z==b^3#C4TGG#g9WPT[84HJ@Z_TK>_eV>b#f)6ESbBNE_aPOSTD,eHg2GL9(#O<]
ZLW7TbdQf^f;D_c_O<1+/3NR;OG^41PB(ea.--Q^ORDd^UB@fDWYBgKG3_Sa_P9A
7=,(0T)K&29S[bYJT,=CB&@E@XSIMV))C@GLWBVJ/<-^4I8LcGTF<8<;VSRY4E]J
fD7?#U[b(LM\<U&;f<d1)@M1a\dC2aRedZD):cIY]FCHT:-7g072=<U.XO008F>8
P0XU&(X8RcS5=BTZ+3KA&N<YMO18_YNb,OA.5OOPR,UK/8M46T&;CIYe+Y#g?WTP
W97G5ZM-JAF=PR1\0@96&V<Y5$
`endprotected
endmodule



