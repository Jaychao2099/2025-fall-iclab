//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2025 ICLAB FALL Course
//   Lab08       : Testbench and Pattern
//   Author      : Ying-Yu (Inyi) Wang
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : v4.0
//   Note : PATTERN w/ CG (cg_en = 0)
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################



module PATTERN
`protected
L<1L)VRdbVUJ)&LKOHPb&Gbf:X:7-eXO6>+D2ZNSf-b[K)d94;PO1)NYGC-@f<L:
A(#ASRgUJ5=&f?4Y][C?S]U;/3NJUUA5Hc6YQD-JG8fZ)@fR:Kcag5b9=_&RQZ(P
P(H\Y\bRLZL/A@5FDD4>9(H6PUB,D(;?e0Z)INT&c9Q_fD5OF^U@)&#fG)>V(W5]
RF5#G3OM\QIUeFVgXDL#4I&Z,b[R9B379a.WTbTQ;^L>B5Ze&UAIcPL1/Ef98A0^
&31/?8.ZF8:+MPZBHQFC:LT?-.ceXT7:+\fQ2d#\3.OTFd)TON2IfYG,0/C?(YM#
cE.;b9/TD@(VJ&L8\+2[9;S(DJ,HGf9@>?1N92O/(NNND(HO#7/]b,\1[fV<IUKQ
J^C-[TN7<<[0C.3GRYD3>==e)L^YZ=fRV<[PG3\\_,7B_c__@I<X9Qc_(P6,H<A+
GL=;-eKb#Q=(-;cIeV93V..f)<<N:YW]<)FJ9L_((0/H@A;FZO_6H[R]UR#CPcRg
I?8E3R,PQ:=YgU]AG3@5[Q6>2_507K2X^,<A5EfAa[3D0PUUbRU[LHLL<]^K23N,
^,J^/&<TNc-=\>AFRK[_Q8&KJ^,fT_UFW>)=a4[]KS.BKT[N>]6eS@;KIBO^I>0^
&V;MeeDF^UN_XM^OO(6f:&C[fQLLf(<BF=B4f4Mc=6R8M-^.Ha[YV[a+R/L)JM9_
ZPaN?Z,/^d:Q5@1;6>U0c/0IBZ&H)X#@T#>R5SVc6J#Wd(5SH.WT]1&Ye.Ie4<Z2
W/H35PaRN=NT\eCIQH[e]\f3VSEg@P:ZB^_=0._Y7M15gc+P>O92fZR/2K)Ma6bA
NO5,2Y>I:.b8&]H7E5LS17CF+I?0g@#HHCB=JOFQY[+D0@adFT#F,FB@JK]PS<UQ
Q],Nd((/S#V0N9DRFF3Q@Q@a@9WZc/7G3W8A6Pf.X9F^-+UJ<VVC(6H(1E1dT+f-
(-+eRKg;c8@.d&Y):@&D+_XS/d#ffKMd7T[8Z(Ig4IaX(;751a7>2//=FQVIE2UH
ZS>JC^_7]Cf&:aJ8;7SD?Fa/[/E<T)&2Z0b75_X939;FY&>Z#Z>C-#,6B&Oe_EON
e?OSOI25>)DK33Wc;7LUJf+)C13-D1bT4+G>TVDb)(Td>0N6@;#^9UW_P/=+),C4
5,g.O2&H?+2T2,J(VV8P0TI:1E7L6(:P01.+8;9eVB0DV@G_;Y=D_<]?7YL_XB)a
^HZ1@?Y>FOM5[X8&NNSBZR8MeE[E->J5G76d:84&;[4ORC-c(2E-cQAVF-bE3aPE
KJ<&3+4MK1S7,gKW?e-87ZE\:Lb<+5gYI2FW;Q-3E,1P_JM];/c/XBWHTX;<(<QC
&@,;LF)ed/C^YI(1cW#3NK=P.L&116HPWWbgcb\<]?9c@N^?#)D7#)X=@0P(,+BS
@;4I4UGc9,OTS;aNTC-+&Q2/)c3D?SZ:/9aZTbe26@<2EJ^dYL6@b1N@>?LK>O=[
a8;T>eQV>d)5;\D>R2(BA1O:fG;U[2Z=aN/3f-5KQHY50H[b:,I22,0SEM6bK&-d
+1/Ha+/\1[F7,&W&OEgEY>]RVFXV[Q6?;T;VWS/JY3(H^)2d52cR96Id.]X4Nf:4
e,3\Vbef]HgdU8bG>A(DM@6c5YbU-ST,6]M/c5;M-RdBV4B(LNMR+V7P<K=d84?K
/@UM=;TU8..2T]4X+D)K#faSMB[]9Y&CNRaI<:Q^H16T-9/2AS9D3S2N8O)CLT-H
gT,)NSIQK1/+Iff_I1M2e/3W5@O88aFD,.;1EK1A\,#VbIV9:f#1#]/9eGIED70D
PZ(4HI.E+81bSP8EMC6#RG9?THGF)a[T([6@ZJK7/)6OD)L_7OeJ]&O=9[1O>M>S
&B2+ASTS6Z[4YX=-HWY\=+]F=][=M4-b),FcH.U743\@H[/D/RNI9aF-2HgS?>8I
\aRL5Q1e[VU5N037:aDABc+THZ;f#HBc(,S6M;cOSHXa)eA8<,W6/?cP4E<?MT+(
THD/R19P&Ua9M]1N5f9\]P[_ce:_cU;5L+QBZL>U:+OC,:E\aV&2fI9XEd0g<FG#
(\GTfFW_@;(_;ag\Ja;c?aCH^BD)J.7:-^Z6:UTT7TX@G)&ITK=gJDHO^2[d.DZ\
TY?+K@D>cCdIJ4@E63#ZX<@:Ug><0Y4aaGd]P/Cge:6BQ2+E[B\Tc?08PSOS)=X4
_QRS@15?7U0G6)6EB[41OV)Z/V=]D_,KY2\)XZR1fCEf(TRX@[c@3af=@G>IU#Y-
Cd6IXb:fP\(S/N5QLbaU:L.@XC&0[>UeeSa6,I(WKURdU-+W2_D0MH+PRW>/D#,-
3-E=<7U_=a,aD_499)^0GgU3^P\<383CaN^ADe19/0ROea/O@Q)3S5=:Y./JgQUE
?X(ADFdH91ZPadQAO7S&K<NH4X:6-c0TM_KH-/8I?X3fa#]gYKRHbI/XE7PHHV]3
Y4>16HWU]cB)-M@F006\#M&]98TaZP1)45dI<#2;Q2eB>(G&9JNYJ_e4/bH/PU\1
9)_P^FAac:&+GL>YMYd[8D@FcXZ,IW6+00KSIIX01(AIMcdB38GF,Z]f]2^/;L7@
.T4D?//U][[_b11?:9&:4Df,+71WB0?e&K.Y:;8M2)(?ZL0FM51B5:T=7/K#X-AX
H(3ePS/UL9,LV/Ea?@bYbCbFaTTB\PDcV7cf1^B_4TK.C2e]8@9;A@0K,.R8cUL6
IJ:)/(3@FB_G5>8@.V2CWb1&a-V.AbTRV8dW+HT;7^ZUFY.K>AEJ[:T9Q^.KReA\
+9Y>)Tb<Dd\D#N)J((#E)+.=T_g^T[>1)5RbG.J3_VMSL4];N8fMT-+Z/_R(BaUQ
SFLD@b,I(<]9aWGO)]gZH6>e)W-Y]W:BU<FQMLY;3Z_<<2+OPG00E2\?,DZ/)@]P
@^G0G:>ESg9cCK3J43)f9)C<TQ>eAH]ND0H)F?S)D[;A?b0.a]:=;5;1D,-Y7LD#
#[V]B+5##CSe&1=-QJ[[-N=PX<P)9.2?:&1//P)YQ0/M>DD,,a9ZY:PRf&#eJ_IZ
&QW\4,aZ:5#P#0:\2(N_a[B;J02&[caEBbF34_-C]LBU#189U/14I+QI#^UVT_,T
3?Q.E#9>2Ga1S6\J;f;6QXa1gM.Pd,58Da3SbTYPOPQJ@H21GAf&186;g]2LT:+f
O)9&Lb(O3+/8CagKD@Z8@#,-Z#2Y_Dc2OR^6[_^H:_U&\eG2V4_WU8B6Fdcg,F13
^F:W?ZS#EX:a]1CI2S5ZUS6<IPI8Ke7AfZaWI51:-&/DgM_V-?B_0Bg2DZUH6;7=
L^B)>R5aM[R(>cJBRg51DfL@W#&F2EN[(OXd<IBUQ8LaTTQ(?M/4Q)=N\8H0<6#-
^Bd5:?fN(Q_bSUUg(f9039I0Q1/UCKEAIJH[G/L=)0PG7.0b[DMQ&0)DC8^7Y>RF
AA?a,3/aP-<<]B15N397TT@A@e03W@]+=VG>@#:^Y(JbSM\^<FRB8bGUJCQaD7?1
6@ZP&4B7gYELT3L=E_>7DVVMNSU=50ON5[FWcACMLT>YOcbCeSCT0>db&QZb@YE0
f;;edEHQAX9BWaDZ3W,T0/MdQa)O&8Pg8G\)-[5+#d+8c,13@g9R]X\BgX/_<+Ja
T>XSaYC+0Od9MgZZFS1])22<BcO[/6>3R8/T<ccZ@aLYKeLGO.M4&\6/0ICK-;;D
;Z,[(2:P22U6O5J:bFY7\Q:ZQ)Z-XV<MVN&=aK5[>:J&GPJ@C8YIUCaQ,c-,CQ->
C2?F576[DX(cN#6>f\(8+^>G9KXC+=1g/9#7@,>&_Y3D<B/2B\KCaBa]R1fV:7GK
6#L48,PY174::aCe:P-6.9S-adO0,57b.]#f[AcBgAA;:5GDPd@TOX?,ZL-KIV<d
@..WSY6a6.7Fc(XPAZI01,c7M^g<>W6?eX1-NIBK9Z87@[[8X=0?<N4KTfSRRHMJ
?\\34B]fAZ&L^K;S/M>6?Je?8AXS<c97>gBBCdN^QEL1(18JQafD\-C&KQ2;cAYM
@[Vf>@KcbO/T#\PdZ#S3e=[L:R9^U]_=XNY>,JJQ]NQ4/^WABM7KgZ>eCY;#KPW2
>/K)6_00?Ue5bG&;_[G8(;)^XV7\T<K=+JPPW5-,L(CQ?9SOLa<-F-7&fGH<b)C(
d4U0S3[a<UY2SJ;=WE?JNJM\I:f0Hc^V@5ec]0@;&.55O,C0Q&cf^=g7.>&HRF@S
-&[W+@_=_bHa,;-a&a)Q7\_M9cMR?@U..Df[)44S1XDG)MgF6@6,)OfD\;BaE)+X
63aO/4GC>fT[eCEc-B>U_7YZLFWZYJ_T,-MR7_;OMK-ETF_=aXG;D[,Q#VS3E3@@
cA+W][Vf]BNSA4U:#37S+Y?fS2C#(GO<\NV[QN2&Z0Vd7QJ<,#7^(NBT#FSP0aH2
DOTZQ=RAI5f3SSUVCJMW20.4GT#:6>Z_2<3?Q_?9fQLa^RG:U8E\F0QM?NCRc@RT
TcN9/-Q0#]U0&C\L]NV^QdF.g+9==JfDV1/W?HBTGWdYdIg5HS<I@H8.g/@/ABLC
ZC70TXD&e@L^3UNQSF.RK?Lb7</RHZC]c6>5RN8c\U]X]g>J8765Q3WK-dd-cL12
I07S<Bc164,e2L4>(d+QKYS.>7TcQNZXJ>X]RY^LFI+H2D7Lf1#c[)7JX@XF>)^A
9JR4_9T0L6b5(+J8GQG3;:+;0f_KE#T+<gf.[D16(B8^1_f;Y,C17c2D/U2bc=C-
59dD794cK6<6b9_5F+[K87F67e&8Hdb6VeB15D6L_B[=[JJ]6cWQX.:fBd&B&?;D
YLc]XdWITbI3;]PO=VI7aeJG_2DKH5Yf:<R2dFJb6\<)Ed^bcFJTR_S,PD^-3YE8
d#:A2gbUXFgX?V_;MOD;H=,?&2D?>ZQ&AZ&g>_T_A?)(>X&Y2FT(4X&b^8;cS6=-
,dHLcB?dTQ<cC9;;WD7SV0GL?2F.b\QGGT:IRfd8F3UB#]P^ONYgQV@W:bLVO&bX
]UDNg6-fPP^4P6@G11])T/dG+SB1c,ZXH9]K(1GKAfN@T8WXO8NB:;K#[(dBW-bR
.[UHA_LRO6GMY0B9K=/KdKaF=<CLI@S&_S=?5f7=QRX_YC:\W@P[KD:TEGCQ;C7U
-VJ>E?4RgZ=cQ930Z(C]<U?f)V>Q],+#S3R.5Y<N\:Ab((6A]eQMZ4,0Xc>L=BNL
NKQ6;)8#-d6LB(NbJ2]Q81;CX[M7F48C7;9@]DK5EC8GV.f60#d=LGH[O<G)T#D1
I?[=82VJ[ZG>ZWEO7+#B<_SB.2fPTgWWORRY5DdU+RHf4F]dZT))(QaU]@4D+9@0
@[-(9DGfR\TTT>cg9&HgLc5>eFYACFO(_T5N5#MKZXLc&Yd[fS9GDE?E4\4D5O=1
4D-]TPJbfL&AHHe=1]=d3=VCN-_@4AQd\bb#gdcM/?^MA76B<0UM./D4>7:SI830
Sg.Z1#)WSWG4?ZI9POMUgYG+:e>9Q.-gU_O\2DgI+:Ye?>1Ef/82I^N[KW2M?K>I
9eUOUJ^[;M1\0O[1:ALPM8]31=gSRMY./fGMOc_a#4UQ=dC:OERQ._WMP<80Z>Bc
McIUR5J<NH83bM^eOO5ZCaUaO0P4-3BW<E4B,]gJQFFNZ_C7]A7]eJZN&\[:85I;
6MLA@bBK2+G=YbLg&6-\[CV6=>D<4JVQM=[UT=-cg50Xg]XgRI<_.b(/<S9N(SF7
9/((UD:WLEZM3e\K[V(/3T5dg.3&VHB+=LT;3B1&^LK.ZVP=EUSYT.]?a>V9g9F\
8[8N^+J7R8);T;B2)YZ,dI7PR6\6Y>\S;,-8dO4D[A0M&PI.6L]cfTD7@F(ZGL4>
SCBMB7CI=<MSN&KY+8fH3[#25O6GYf:?7RUB1He+MXB?H#O&NYdNfKc+P.;DHX6O
PN;G:[N/W1K^g5P&HDKaTJ(:K5#D.9CdaK^XMJ#L50aRM_J985YaFbLb]_4RSMH+
FSDY9[&2)1L5af815f2-,&27A\&C5,(D.4eDPEgaFGBIc(KV(cX,U+RA;@?T4&3#
V7fK<#<cCO0F:aQ_+E[]>dJTQbXYWLIJ<9=+Ia,<:+-RS[N?I9>_Xe&[^/V<-UOU
L9IVcVddKS[+M<EO\5T:N\;e7S/@5__^aB9Uf>^R^&c98,GR:OF,(9.23:O=]I6X
6/a3-:;@Ub+b&ebHS\0I@M,b5W21d_KZQ<C-gTK\V]#Y/XJ_CAb5I;TTLX=D>_Y2
FN(BcL]B?(bYVN[=MRGSdN8S-DLS2J=58,eaE4XM-T+6KWMKa\56:C8=J(g3Re99
a_AB3P&N\,QB@d)d>]Lb_dEV))XF#XLa:.92R?Y_Oa#NHC44:NUF0a@[[TAH>908
&YgAFPF4?>@A\#;d=dY(W&X3a&#?5NCMF3AE@B/_E86dYe6(AC>e6AI2K,0Q+?3f
DG^,7g)ZNNb^dW.PZ0f[2c&gdU;Q4RETbHDS>Bd/cYS6?W1=aX(1](I78+C4I<.,
d)TdGa[)8Rc)5\bHgBGX0F.2=E5^WS<Qg_MPc5K.ZJTHgd,f3C#ec8:U0fFcJ0?8
aH9&a:I07UKdDdG91gg)Pa]@9J86J-8f43f&VC<OM+b(b9&E(^\P+;<dRMV=7)0E
W3=-@g85?1La]<C\7..YEI@O#Wg-HS]Z3^a[X?Z@,VOaM</bcFF(Nc;L6P<62/B9
#^UTUFS@QN<,;RgB8<U+Db8ZaP;+d#[S?+FOJ<XA)_3TPGZ-9T#DFC3RWPZNPFcL
11e-G6Zb6O[Z.J@ab3&O.K^2P:7.-QCP+=5@(LW#B8&OQ_bTDC@NQ3@+Y^DZ)Q<J
];U&#KE+7c0,VNVR,dBO@=+gYS,3VM^()VeW(CaWP4,V^/H[LHX^/dS;9-_@OMaD
C.4K/&=SWYaB/3Z&eHMTFYTBeENA03c#(e7e&5<F/.&g;=7I9>Yc1PdO_STf[5-/
NZ,RK]Dd[?2HPJ&aKXc6X4dL;D4Le(T8FZDe#gP/5dIf1P5f4K7E_0O0=8CANW+;
0ICV1ce54B.Ofe4&_e(gN/,fCW@5;?-d_W5g(_R7bOCfOT\YaKNJ\R6F\\J4_PU,
_3+NfYHGD_\?T=OG;5.:)LB>WHG?\g5e?AA(Y.A9I9;O_Ue.IK^,]HN)I,##N^=F
SI6/^gOQQ-Egb=_ea#34+4D9X;b0NSP3S1b3HCT/ZNQ[3_L733R/8GO]=V18b[3#
U@gW?M\(URHVZW3&2\)OS?1>]UdA9MS1ZVHLS__]A8eRY_YK\-<cR#bGS&B;g^8^
?_\K-M?#)=@)G:&X/[371-OPG_9a6_3/0@1CU;SeH5dL?BNfZ+B)a4=W[=b\[X@L
]5/[>;54)AE9^R1DeYdd:_MQG3=5)=Q2L\V,4.04:\R--)+?78fSVII,a\U;CAN8
J]H1E+ZM8?8;\)8g_NgUV.VGAHL,\=1N83^^OU:<VfTaE5;a&]G18ae7NT0eMSOJ
)V:6/3HNMb2WSF+Z+-.^bQG?3aKO150Z61[\/._2b#+G[[\&JQXg08UHEC0&-&LE
9fC@IL2Z)B8R-a;]dRSF6[g@J,#e==gKOLcK7\&efA-NP@>O&\YHCUY..?9MdW-7
+NI2f:_We)=.b4[_1eaH3V>HPg7,RYf:D3TB?Ng.ZDPT+HW^L4VbGI0#_Hcd@c?1
]c\0?:7_]_@:<LM=>08LDWQ9S6a2#c[;]86G]]<RTG,@1G\4Q4,-J2LT6\5]D&4g
dDP2;<NT0_\dP4T4Rd^X/R>(GI&2+OcF8ZCa-7)OA=J3UgTLWI2-ZO7d]N&J#5ZY
SSI/X2-=M3[=R1(S&]-XQNH>@>-Og\A,L_Z(JYbUM]W].>F2NQRJMeN9\9;/eB81
e\8-#.F]X\7/DJX]a[^?MVNZ:&AY?NEMYFYZBKC-0a^Y_VYOUY(+?OGWC/U8N9\a
8TSYE^=ObXJP5C:R&;0>MeV?I1:Z8A17R9M6R)1]+K&E\T7S0De)IUSW0TD>,gH8
BXD_ZZ7,8Q,<7R+<C&(CA)?65<P0X#&?N/bRYT=Jf1O,)2TA+7]D-?KAKP:M0SU<
C#QGH5G^8IPeU>(d]LT>FRLE1VCU+dO#P>;CY@1RFeO],/7Qd0=MW(/Z;XZ]C:V<
7GeAOM4bG,ePV?OCXRHf=2Lc4JGJ_;M?;^B+1OW,4BKH?02<;;1G=42?0D/NV\WL
OZQWb^MB:AfR3YfP\dMWeVbB8T@V/JB:KS5QO\T7#)SV>D86]4-(KYD:F9<7([56
cE<,G6N6.[9YCMK3bK580^HXF/ZcX48GU#e?SYd:+0abOX<0&(UNJUPZCaZ1UPde
A4af&,^K:(F:dg3EN;</TRGT^U[]Je]4K69]3Ka.d^,cVAZV=9J:68)5B:4P46>/
DN^<H4[?@B:e-YO6d>RA_FPP4eNQYW_gF#1B.a::O1GC6@Oc1dd)@8LOKaY1S_/M
YYJ\V@aMT@H.?g:D^QQH5#XSRS^DUDJS7M<IH3]>d/3<)6a_IXgBg\9T6JS7]].V
.BNRP,Me[B^8P^T^2I-N04GXJP>d1#@AEME.VIcS_cHP:=@R[U1TZ-#NfQ__SJFZ
cK@c3T8:(bVAR4WX8:E@85Y?PgH)&O)agU73-W-eBd1CJ,2g8TOCeb9[,[56Fa)R
A_0R(e-CW4bM_<IRd_Df^3QWP4GO7I-U&F])QV9e-2d5]>e+,=B,4<A>NZ01gL1G
2K-+A2T68R,P-8e[?G;3&:F[L#_,7cc<JQ>8UgLef54N&-P#d2bC>6/9&D1)L\CE
96O?1;S#\>DOL:a[Od\32P(e)16)&P^;1[><9-8IL8ab_/BR3Za7d),Y8;U\;A1E
cWc,[88_.SMCUKcN]A[>I-9PCNX)HA.A\.NZB9CLJG8Z8N[@T1-0R7J)9K][_UE]
#@DZ^9Q3AZO@a;>X3DR-2N=:4+Q0]B7aeY-6;#d+:MCY4&6FWRESBIgFR?8>7K;,
85g?\dIKLW8AT+5cRYg5>fOV:\gJ.C7(Ve,g8aY[\8IcA7I<9Pa4(cPJ[/?(\R#g
B-F;S-IT8AK57A885L,3./fd[gcP^@N^fY1ICY5VJE>MR)]X>:S,c#EJV7A)N87M
++9gD4O^fV]U#.SaBe9H\IC\I8?;gCU<6J-#<ZQ=OKg^<L-LZ>09X7G-TKG>#)?8
R4M?DDeD>;C_D7+ZbVCaW\=M1g-c4RUN.0@5#7^Z]PI^01_a/7J4#)4GYT6JBR(;
91X_R:@(9#/eBM\?dfHQD8:T@Vgf?+\QXeW(-9EW1G#WF=44/_Q(KEGLC?5MN@>X
eT(W2-7^2E<[]_[OQ/4^^03CcS?&>:9-(8QW5&c@3[T_YG[g0a&9]gO]SfRDba/2
\F?]C#4.VD\GS6;Y,+=U.3eC6IgU.?=X\4#EZa0S8:fFKd^3EI,e>]F5>13K2QYC
bad;4PWg3N:-/GZV1=)94P-:F,2)]fGA^#<@9#Z<B<]>;H]],OVL3a8:fMIYJ_^[
(RWBL(e5V,AX:]^K61EX;6#2X?Y<JRQe@\UK/>daU=]8YWK4<;?\1aW49aJO(fHd
4Z).-)_9>#=TTDc(MaQY75PFV-cJ=.UaT)R31fHO#Q+6[QNQ=gO^=>NSWd_?O=>L
3;3:/S]2Jca^ZA?H-HXb7W>#c;)8e[eZ/<@]cGYN##/b8)W53IOE)Z<?4NZF5L@_
8I.3C1F,;bf7QOd(QM6FOK[:MTV:)_b#c[(4C=eb&=6JfZC,5]d.EbON/8#>f[GO
=G+eOWBg8bZU#J?@IB2/W6[?&\V5IGfB<V0fK^c(d9J.^AV[:#X[U6#ZKg_HHZd[
dDJ/2)>CRdA#VbNcUT)T9U,CM9dRFff\P-FU0K63H?+/NW9a03V7]0@(G6JB?R/+
W]d\6,DgBR-4PJ5-=-a7&&:JAL>@EdJeY(Q)GC+]^XGI.-CW=Tg,^<L&?CCM[IG)
<]5PTX&bGPA;Q]PJ&2V1Y;(K>PSVQU\NGY8K&/TP24LHNeYL^bXE:e:I3HOC?EX=
/=30,a97_Ugb=BH>>AJKaBaAe_8_,(0Z+T&>?J#R\;f?X2Be(aV\WfLXZ_.C0_0N
RW@EBV&,^P<)L>]H+8623d-Rc.K-N2<O9>GgVGB8FdeM]eN02eA,TR+T=9X3MGYN
(I]fKCVLR+M(GJX68X(a>ZBIggRG+ZE)&>G.;DD,LG.PN=1_<E]Wd+cP7CQVbTE<
PYXNQPY8?,8UWOP@Z1>7:D1bPAXY;NeZYPS7:GJ.W).WWQD0;DT&G\@<b4SA)\[Q
I5IccVf=fP4UdMZYgO(H@W]&,g6TS<G6:.Z0e:Y53ed@g5E.71]PY5XOGY/faYJA
)2;bG;I_DF>4RB\->G_A@/;7QbW_8+D12D>K/P4D&:=U;5;bf<#)WW^LN):SY,JV
+PH(b1Sgb1]_:4QG^dIQ-b;T)&-SYI;+7TL3Fe/E:bfN^c/f)K.<2MJK7PZ@R]0T
:<G3XI6bM5(Nf\?(HK:08:BCRbA]EA1DR?YCW2<CKg51]Sd)]6&_4_OUBS\)=Hg:
4DY^_M;-D.<b\b;PVU0#EIg(^V@c[/6.^HAafg-S\a^(Nc9Y^:A2III&R/F#D/:N
#0:<J(V;fH.\f\Q(Q_GXZZ?S(74_DB?Sde]dd:A-F,\Z<7e<#21TTL50FfAe7VJd
22,9IXXU-H\GE>dW>+Od<H51M]H.T^A^E7(48QM15V_CO63;XC=INdW^>9\G1,Ed
<WA5S/X^#g,;)-N[0(]TZ_ND6AHgcH@U.OAE,faZ&8>LCAZ]@7O[7A#5U8Z4R3KT
X\)ggJ.LP4C[:39KWOcJR2\T/Q^:EBM^1#[]b)MEV(W_W;^+=U]&fT3O8LBg=NX.
2L=fK(GgM2@EcP46EEJO/XSL?CM>+7/DITK_3Q_GX8G=ZgHRSDUS7fRTO>85I7e6
dcdTLa<.4B]R=(G7N(>.,Z7YFQACOO7Y&G/C>eIScW\E29W>1c(:HVFcR4fL&G^+
&1Kd>AGQ/<9PWIBW+^B#:+daFFXX4EI?AdL_a/D4#_6,]4JSS]/<b&/(#EU)-Df9
14GaY9X[XdRa^BH;Fe<Te>3U6^-U8WB:#]W6H31A=VF^1>9F5:&^QX@bc\WCR<Rd
/FO_FW/)B4)R/Z==#/[eg=I>:BMgZHTOSQE6;XW1]ZU>,YUYG5fHPPO[-X#f=9fO
E3(8g9(]@T=FV\3e1D4__edND6OW-QS::C5L@)/AgMdLL^N@;RFHeR2:/4AX.bSL
=-bJUe8U/M&[aI^WYI,WJ?7b:0#TM_<gN;>)-UJA\<3B@Q7V<K@a\:FJeV4^WUC)
3S[117/[4+8]1[N6a8A+;P_:H(cY5a.Kb4GSZPL-X[I=I=Mf1g?]GdIYRd(^A:#:
#C19]=]ggAcUfF&GO?(4+\QXO]<VR[-RbZG.^M>RL1FF1@YPD/SY(2aCb[da.F[^
,3)SDR?.].-eD4_+G(00@[?6c3XNGZ<COL<O8cE&-]cA#(^NV.7\ZZ0Y<Ac^4VaF
H8KLCUIZG;=^70c^CO-CQ\H;:1J//.#FbS&g<Og,KG.,GWX[:F6MeRfM@dgW_<?d
MB(4-SbdX2IKT]3]:3;gV\;^30TA106Y3/(ZY1R[>_?Q9?_]?YcGZTd?BS@b#dad
)Q>Mf9+PCA.PZeEI^FP/e&Z;?XE@5+_fcb40A-311J(F<DU[9g-?e3gHY]8&JMQ?
,X8XX>-R&&4g+,#8?XC<.8U-KPQ[;D96S+,\bZ(/:>@;3#M79[90R&(=<144fB=;
^J_V<Ic@6aaTM/J(0.-a<8/:I#Q3Tf1c(@VPSFX-?+VJ\bOV5;DF2^4=XEg&d9=_
<DBfC<1<(VE&0NO#1.ME(_8YW\@P+I50KL?1O_R@g_ZSC.U0KfTEGcY0(V+(_MJD
E:_H;IL&L^c-_&KZ6)_;gRI@M70UO_LH6#gM_78#2c_@1XY?\H<UFd_+5E)KAM/G
X)@-3,+AK.+dT&fZ+XY<V@B:H&EJ9Z_@-1>.@2.:2WS5^C(0)HI@8S/CM&(Q>)8<
)0^^2C#Q/&6HObK]C&0;;2V)GfJTRY5;R0Q@)#.(IJRg-4^&)=[LMALN,62]-#g\
>&8cR:E++QgIEDCc+b;:/W]SPHMb(;-FWNC778D/4cA.;UL?cN9VJbU2+^XeD/L2
<G;RJDR>Ae3dG7d#3_(fUD98(+aR-)DB\R?P/7.R0Z9I4cW_,e1@PN8Fe0946K/4
@.#b[3;E9<.]H+/D/<T+D70_G,E^7(2R/?@/:O-YJH:AbGG>(C>^T\e680ZINJK5
R?:#[BRVe6G64,bP7+][MB/<b#O4-]D/XZWCIC7b;:+WJeeW10?O9/9J(;-^TBD-
&Z+2RV1WdIH^7.XHc1HNbEaQRAZFf_?_K_S)7.e;_,@J7V.KdLCb++ePPVJ7?+PZ
;NO?&4U7[[<SNB7<SV4_B2<Pee6f2Pc+dNUT\]c&K1RVf;5^:8(8YNFQ+QLU-HaQ
;5^#^QPJ(F6NI&FZD,T_8>VKcW+/Gdd/Jb[Y0W5/b;cfbJ[+Ne7C5XTVUdM]X.][
3EJ^,/XH7NWL+[,=N.+5RNV2\=WK^/(R?NIe?2:78U>UW#RHL&b)8@Y6IL<JK-B0
D6ARNfJP.U3YSM]Yfd7W+EHgGV^\<IZc2N)UOXFKS.)7XC2BW2LJ9/GLTT-CE2WA
(O3O15&9Z?6G:f+W?>PO8ZNN.PQ<P+_POe,D_gc5+4AM0#4@a\7\@;8/U)7O3P)_
fZ;XD\<4.N/eW9<=+(6@\IIZ:IbBd=QcJ)HaI[8IB)RMG4=,2X.YJ&74E+@cC,R(
C1+U+S_EPZ[]f2:?71.#P_]LCHOX4H8\N@SJ6\TFg4fgJKfb9Q9.7d5GEEF9A/A4
\:e1(4TG7Z>H)L,1aZ1d9?AEee:(Ja,,(QIARP&C7[.#2=0G)8WE)O^2:@JB\9Mg
b1KD@c@ZJ:?gN:A@E26a<A2XXG,SV_E-X6;gSAX+gU[C0AWb)&Ec>9?[)b]CDD-A
X8.,I]\fYdZ23[bd+gK@#N<H>3M:ZY?cJa^39PBQ@?Ib4Sf0d/P,E/I?>LO5eQ&S
DV6]<#8C<&GZP=4U_\dcH13?Z-6UD3^Oc#ASOH13eA<0Cb<++@Ob]B=4I,8#,Q#(
-GEfc&419?5>>_d=H)Eb;Bb^I/cZe.9gUf94.L29IWGVVWaQWaS/)RG_?(1)[Sf+
RQ0AfZ#XS6.fY9HTL#B=##48D7?0(KM---8E_25[J?_;OZ/YHJ+8^4@C.&ag<I^R
R7FK6-U:\#8CWJ)fM727JOA0;.U6+5Sc.4dU@38E=e+#b,^F8G2Q>Beg&_-cSYNg
4,],66Y_N5+>a<2VO9RU)I/1D&5\.ILYV@NDOM6aLdDN,@)384@FaF_F<g?.Xe/I
,cSKNL[XF>B:fC7)8Q^e6UIFWC8SCWZ=I.44T342dad?:<J\&-G663Zae74G2V3R
=D#A8(M4I+A?G4>fKH&fBRXSgXS?IH07X4&=b:Hd7.04@6a:9W08+/NLaIKY,]N3
WdL5LeNJLARI\X@Bb867Hd1A6>1EPgH:bd,\abRb#G(?<(gJFXO0Tf\WYC1C>4R-
]^TJU)>?[&^F>DZXR;;C39_1C.6M]Qf9].RUL\5(61_V-<)I1[JHCBS?=ME&&0DM
N2+MLfFAHI[S;cDW/#dSAJ\g65Sb<YMNec5&P,3\1Xf+Jb#/d+@+)]IcRUeV2R(8
DSO?@d1ZLGE.g+338^a:g^e;d2,Z:P[cY/CAXWTI#C49@1HU2&<_6d-gJ>5YfFP_
JQR46J,1QX=bcG+Tg>\4?,D3gRXOg::3[;\S4>A9,WSEa?,(::<C>-b06<TbGbaC
O#8<e+)HISZM1LNdD2B:Bc]([09WYFS2;,&8g/WeST<[8EW@\D8]DCI)6?cdcfS_
EJDVaKWS6849,;\,^d2+;Tf(+>@WXLGN;U9gcUA/YB>f141H?gd)+_0\IbF+1G<B
^_0@cY[72[B73/\V50R52K^0)=<a0Z_S]^O,(e1KTGGR<6GEJZGbBW+7[f9Hc6RD
@7[e5baWSc0R+/DRQ\a:fZ)H64J(e))\?XC;ga;HS0Y\\(TQ/SZ8.VQY\2O_IZUc
:DJF]^g5JR^W]IE?[C<g:dLUQb^K?.#62F?^g8^BVcM.T<ZSMeDcKHdV/)=</)J.
I[\QBNEY;A75=+)QO:U/R?9-4;E^XD-\JEZL/^4B_INf30@#0fX(LS[&84PM2AMe
MKE268TI(=Y.+P892<W4X90S6DP(dKQ>?Pa.&QUdRe;6&d9aFF-MF(aIJ8de^1UK
\M;(>UPQZ5GNLXgQ(c-TMD05OE1,/Q0JSWf:G?7&>EE\8IW5Ud=COY4M,ES?:/;g
V@3=7^M>7&8Q:U[NUEb,=CD(=1N4(\^FXD)dZg\6@D)X6Va5#6TDBcCdX7L1P[I4
Y-c/^_KeBAEA4I[E;WWMHX72aYaN+;^<)8>CL]gYMG)1f>G^?=:76@f.G7d6R2]3
MQX58#Zg-g\80WD_2-?V&0.FQ7PF?X#Qb1+T]1[Z5HLgM?PP#AcU7:IaMAL>^@BL
R&,E@=H_[EMN_QWK5+HNM)7@=gOC<^55^=6M=B]Z=Z#TR7]TE<DE75LOE]G]0g:D
DWBI6O#E+[M9.&Q;/\UGFL8WPF&P>YeW@9>1C&AaMObcOZ3W(&.:RHdgF5^EXe\L
bg#/&H_JIeR\=3W=NER5<A175gE@_f#Z(aTc)d9K@9J2G1,;N2.QS+O/9R71-Da,
fY^AWGHbW\I8da0=d0M2EB,4=R.RQT(2a)RLg)9#B;,6bG)a231O59@FW<K<?T6W
CG_+\/b3<1N=3ec-FFZ_]#]9(RY^/e#6=,AXV3(O;^/\99J>=1MFIBQ(=O3.[+&J
4e]+]+5-UM,3,QW]bV@9G^XOM=>B>/.8d67@,Y(-H<J9cK4L;C\<<:2C)>c.5+<;
--?cV(QY)77@3be):YdEKJN=#FefgObJg5Z.bTUD(X(A,+aE3HEK+3T)CS1GRgTe
F)#e#H,dMdM])N^I3=e&TW\JO9DQ;:0:T++g0R#gVRUN>W2@A3?_.CQ7#O1.-W4f
aRO4&eR@=6@?Q]K/Y.99_gB#a6eE72ZA@SWQfc54D9?3&@&.<NWL-f-_F>0\d6XI
M.AZc8G2L(X2?)[2MZSJb8N:-(5Fd45?aJfe_C)(C(>:/Hd,GN1]f?#E7b:RGNH=
+BHAJGR6-FA(\,,R:5W_1G;UO@b\OdJIAPLZB,73FWP,RX/XW=\0C^?PD84T<&0g
V2WM@>,YWAQTYgKTP=JXf8SU+HL8K,KIeYab9^1=5XH,[XJJ,]+;H@SE0C?0:)_L
gH>YUF>Of)gAS_eGP1geL]3,Y7C@TLPU.,;Y\dCE+B6.FOUN\O7S<H,VSA==#7#:
D?\S[G/[HgZ=\L.GbU&/=d\[>:U:FfN&UE.9)JAWHb,1@,:KTNCX,bAWQP1X+<8d
N-.gVB6@33BB86@[b50J,^-Xd=TS(RDc>L&dBe\D#Z+-BfKZAdB#O9QRc@.U[3]G
-:W^J5+9KCYEYNQ982)R]Y=HCbQ&3D4R;7<4?@KgVB_XHc9?I_D;?#_)TU@Hf&<3
PK_8)\2b(]F[RN.0S35_Ac)O2<8Yge_MH=Pe@7,g#9gaXc(Pa6KH?_DF14)<<68^
G5J(6cBC9b7V@C\>S?=;KFL+LCCJ#K.LCFFe&-:D:VTCI0C9EaHMLXBdHKIPJAE@
TGS.HQ2>E-fd/_]<2SH?Bf>6^-fDgJO<(F+;cf)KWK9A>Eg)?&]0<af@=&-I7T:1
YC/^+Z=0R:34+N+Qa_&=P&SF.[\F;LL72=5ZIE2LF>#cZ3<_fgXWb\SPH=JG)FaC
+2WZ.5YO.27b_HY.)3[Y1NI@0Y+bON5@M,ULU:#;^8KIbWFDV97FZELSA3f6CAb3
F2CRS./W/SZbR;SS_45#Sa:.T#@+NKSC]DN;?Q&O3FKD9MJ:;I/;Q&;(e_Vg&W_C
]e9,0RJ(7\#X<:JE,5IC,_09Oe>,]YY&MDUTK+KNc=&AJAQR(V&KMF67&aHRROA;
\:_&X)./_QD2C\=:eLM#TNVbTA+)OYO<J+4)eK52[@5b0#-.GN2.0-N&6KVK6C#@
=6.B(a>H[<KBC[HAKEA?177:L.YOaf)d^a4A/Q.V-Z60>-Ud@99d+8(<@7UN>MHe
bIPa9(F7IN;a^7[Q=KY,(?^=caH7\ZHO=+O4^A<+c&2Be=BJ-/W[C&-6B<4MKWJe
WB-^Zd?.P#_CDBJC-^^;2]\>D?Ra4-#=>+PX8>=ABHD+UTE>:aAYMR9_=MSA5cTO
5?EIOAM?dI=@M/I[H,5H1T\;d1=/=;YW_0BOe^3U5+3HEObW+\J1<SN>TJ6;N=KR
-<DA#87KV/77+Ba];9a953QC/?eK)80]8@af+_4RgK[3X=K.7Y;35-?69IK>BA\d
D6DV]VE=PNKfYR?>OM>U4VAfc,OZMdcX;J51<[VPN</GW1+)Y2>O8d^GQM^e\G2U
?Mg./BMG=CP,D]_Ac2OMG/G<1VXO[D3ee-GJ(Y)MB=_f0&4>-<:GgPBO)6^e@PAQ
AK1;_C<gI#K(EK?8F)F2?=Z?E8\1XFBUKB-7UME?4ba4<EfN_A3/)Y3(ZI^K/WLZ
&f)d@?EY\V\AOA#g0=IcE+I-J&:,:[_(f&WP^K<>WB(B@0b18a#L\LXHF?-_7628
29O/S-T#V/)925cd_aCQIc4HEY+\[F7UDFPdO4S0dcW:>(M]GTY(a\S/[L@N.?FR
?LfPCMF+D>>ZNWLVXPbZW=A3H&\ZB_HHEN4<VPBQ?3K+fb7\d8<IG69e>R=RXLYU
K#[9)XJgeH\&/HMG^ad#^]^=6D(NF)e,e@Q,-7;1AR&T8Ka]8,@YAE>ZEW-ILTYB
/Z&ZC6AVRE\1S<_@fXI]DMYW:FBfZ3[0-,>F=6)?83K.S0f6-R4Vc?2PW5;7--29
E82&LZ.IE?Q\X[BP.7.?7\U-W=LF7.dL9O,97R>8T7-a+]L)(YXJ_-Vc0?OEBeO+
Z/=-F@_XT)XQ/T>6=^_Z.Yb3@5BT#,-3OQAc9e=bcKZWF.7;TTNVeF:;YJedS13<
DQL3JSC.-_Rb\57NJQUB\Q6+R1M;I/#0/Q?K+QQZOSNJJU6^4:M4K<D<8g/YO@_X
R.BUgU641;9:P#)1JaeAgDJ_7<J)?]D4.cNS/c1)A:6a-/WIZHDI?15PN,--T&8S
5D#R;L]))P@97_B+\3_4Gf-a7C#NKS=9(LA-&/Z/\;(C@HB7OEA^5d8bF46=L]:Y
;[@=X5841(WN^;;-gTFUTUG4/WT?1[2e.^8b#1TL9fL0KP]IA,6b5a32gB]4A?/Y
?3FdN]3cI(2\HP]K0NPZ)[:OZ.QJIW+VC,4@d_J_[FP:8&E_+dB1BSf-;Sg]I:7O
)O\2A)C:]03,)dQC)(+f)FGb^a7>De-JO^5W+/],Mc9X),0QED-M+[SG5E<\>,J_
9bd4M0cKb,Q-<aMZ-^aAI\7^#@ZScC>fO:6<K#>Q.;:W8Y8C:d2Z8[.(0dF]#[JH
CR/C?[7Z7O#WDVAP8E4P^;H\H:,b:4<&VOG8;gYALcI#NTL@H)UJD(B/+_,&Z5_:
\N2:0V2\Q-6Pd6dN5BBJ4:LP14KdL/T<7_eS_;H0a?g_.Z+EB+,X9\FV5F>1?,.T
384YcIJNS41-101<J,fC8:QGT5]3bUM:Y0-Q0B>bH]fge/SU@TJRX.<JF/J-]\<a
_U=_9H@B+P@JMS\JMZ/6A-4.<?9+L#6f>RA#H;7TP@ZJ7Wfcc9MR9-HP6DefQS\I
fB9gT]SE(F[cY3U;A?d,][@F,I5GMJd/5A,8F16ZD-@;[P]JO]7?ccGZ-T@FD7R5
\\<<GVQcPH(]E?KXEP:6#:_22NaC<ATFWGYYdH;P7:[F#)>@];QJc8DE/KQQHcJW
7\2W#B<L<,8W[,5+gGZY@LT,1^4+d/NE;Z[MUHDSQCe@D[._BPXD?;8bOWb.&ZdM
97ef,16f0aA)Y8<;W^YLdaNA,64a0PVP/7;:=BNAXW>P?cN92-V6>TCWAf6N->3e
1IeH,YJ2F<c>P,30X^YSC_STCM7Z\CK(6@dZ2CgUa&gM9Z>;eU_#[F;_57RZg+TT
CR=?Y^R;O=XHN9.>Bad.<3(LB]aN6\d+9NRbTX2a2\G^8SRN1bcCI\N:[YaO13EO
f04&^;H^ZD-aa7^gW>dfZL^+CBe3108J0K8:YNN.RTLg\6Y>T3(\P5OG8S7cYa.P
Ye4F;d.YR,Dc@1f0@D:+<aD=RYW;ON^bCXHZOA&b>@ALIefBTC)HRCf@e=<8XV&J
UZB?PCP;gYg+>77L(NGWD87(3<B<-&+,fO:P/_CF#e[aOOe:HGFX]N]T/:YH[fS3
Z_:UgYScGXd9FH-?_U,MaJ@c=[BF1,\YV<469@Ze._HCQ:gK9_.0?G2TN\H+VHY<
cYS.E;J-e46-^O1C8W[\V>g_DEQ@e17EIe=7_W]Y47c?QR2:7610a7K@F:3:UZaU
J7#C1HHI>U3g8,/.YXWRGG96J.P5O,H3-SN#/aVOF,BY\-:[M7Yd>Q4K5+dP39Kc
/,&,Xb719J^8JbPKER(X<AIbD4&5N8g1f/]T<VNc;&U,<eN3PRQdaAJ<ZO,6ag)X
??AC;G(C3R&U0.,9A#F<DG)DcJba#fbZ3FJ[NYaL??@?YL0Z/E4W[<PN6GYKX-W#
b.].WNQHT5F-,&gBQ(DK5HD(L4cc?8a70QQF_>P5.a2fJTV-,&b]a/(Ufc[A6<L[
(L.4dOGg,C:VRTVR6&d;+B143#<c[1HRg?D0KZ@L_CC2=HAYcJZLEdB(B4_fX@O\
:HIAY]ed[(/;H;F<DOXR#g)gVDb_LRPFYFIL#;Bf4C@\fY4NLH.[aSE@GE=@;Z)3
Q,[0FS4YV:?SQd8a(,dL0LU;5_P2(FeY6QF1d>B@QOB^)0D1S.9_R-f)@,/C+X:O
/+Pa[K?1W-Lf5aN\dVJC+FZ/E0e[HcXb1d+N]NJBHP6.^3@NPNF&F5?-5#f8>aKW
UP/<d^<_)_0g^[GB.?:/YWRWHO=RY7H4?O[DO:]dS9,40=Q.g39-VMfM1JY;>@.O
<4I+S7J&?B.>#eNHL@OHaf].[=c@&.4,f.U(FUD014\?Q?M<ZaCNY5US^3UJQ5+e
A0#FEW)]W8^HU-?>P1bZHK@7^;RN)8\377W:GU[T7=Cd83SPdXG,,N>D&R<3,LZ-
/5;>F[[80Xb8?08DA6LD^&>+.a]25,1g<12aCEPM#=#AG9PBePefR9^ZY9F;]845
A/VXOVGYKXQGI,eK)H,1UOA@Vca3^fM]_g8P,OY(K&,&ZeRP^^1S6/#f(V/KHaU7
WXKW<(K+>B0M2#@KIBJ.WL=7bYP,31&KJ)JaQL4/:]<T?2HSZ+gOK=6e?09,NX:d
8aX08JQ3L.)G#0OFd?;9^dXCNLD^]b/>Z6bE3c>OQFI+053)@PIXC:P<Y=3;UH>a
GZ#,W<,VS4OU8:&?@f,VdI2L6QL/d+>?UU)(?E<ZOFa]HIaBUQK7d_)BOeJ1ZVe@
a[&3<HUKG18cSF5(MI16=AN^IN3gLM=T9BY./<Ha_I4:#fKcL]IR4I=,B7e-QUb-
9T+JQ<2f7,:/>a-46.BR07B:VU#F2T#+M_O6I+aTbFC3JV18C1N/315ac#Bf(dd7
FOHeG8)5<TN@3DLTO3<086c#@79RIKSL4#3][0&_M1#6S>U[^DDE086e]B<Y+C4J
^W2<+DWT/+\Q&W/dX[V[LWb0cf5X#7)LIca>cCR6>gF?ZcJ:=:+7d9HYK+_2WcN4
_HD_^->JGOR9AL&VP.EN0#/N?YD_?b:Nf8<L^S@R3X5Z2;M86f#b<H1c+8IB5A30
;RKEg29f#bA;E),ZTWF(_LJ-DP+:+&H8LU2\[S^E_WCD:1dTAF8,cb#6H>@8]Z<S
>SQ/(0R=G;f>)L=S/)?#>2OU/_7CG@D/C8]CLO18Y3Z0,,cUSd#ZNDcVU9Y[@>=@
_Ka\Lg/#^)[@bcBI/Ne@>V/g#R;)Y\67>DMJKX0:Z9a>8bW?+KR(MbZ?:2Jc#7dL
;R1<Q>P&NDc_497L^gX[AY>bZNQWU&_7B0SM?bJHbDF2M-9SOcG4+JJ6GdO=7(Q-
V<V)4/26E2[Vc7JVUI?N@aC,?57)3VSMZ4U78QFG<aRH^0Z3T9cGW93>BXdHVcbI
=FU12bg+&MQeX)H^<PHK7Wf:T^#Q5_bOQ7dR>d)?M>[D[UE&J9f85[N-2&VS;cd)
-B8?+C7\g9Q&8a#R3Sb]:d,G#++@PYOW9ORH0UJUOZ(RV_WV6?CL21:;+AffK68W
M<8+NR,;3@G;ce2OO/1D9?E^3Lg6\e+Ce3eA#U4.[BU6,6bZeI.\D:;.[,0EG.68
.7=03762S\<?(-@II0Sc#F8NH_eQ7GE4,F/8CS+F(MBCdS[?\3ZLO<]CfQVQf)]=
E.UgNUPT4DQ.6AgdJ;XX7eE:UV-3UX+5ca5#UH>A2b^gf@F61fb+_.\;>E-PH=M\
3ZPWgW]8UN>;?42A#9D8?L/+YV8:H=+bP_X/7D5ZFC1NEgIR0/Y[=#?ReYg4CaP]
WAMGE_0(=I>IPCC7]<:Y-(e]9+ONE:JIX9[<JHRVcf/=b[2IR\Q@Cd+/0BC)f7U]
OA4&c@4;<MPa_^6E[TE?^23#4dccG4[>5c#Z_3LG9OO=O<G5/bJfE/[N:9>U+E-H
7c5>LW>_84#8XJ:&b;/4K94<>C8U-(139)6_S;(Ae)3H:G1ONL@VaBcZXTJG)4XW
@g=,YI.2C&3Ae;1R^R(L&#G_HKPE]B^DFcY_UTZ/=/J(5NU[)A])2Z5QD83[Zbc5
Z4g_;C;/ND>J\6S2^]8L]0-+F8CM7TDL1W=HC69H/):PLKG3.U>FB>Q=^Q;_T6P<
YX\5E+9Z1M4/H]W@-NZXYbJFXG+2_P,66/&X^C9D@1V4@-fZS+#_ZZZ_aU1?-<&5
L?1W>P:0I:?d/4K=+[^T1\+a=Vf@X(/O#(8Y\Q(_22JK[V/,U4Z]/B>KH,.gPf6c
HYL>M#B/VWPN?8JA/IHKK[41;MMa.Y7aOOSMS.,4Dd&6;E7Ad9UK9K7K(f^^Y+M4
X3dC2(G]>g9T:;DQEY2:C)b5(LU.fc0(A/5SA_aE>Sf:S(3O.;g9f8U_cE#_SM:9
CO.XIOSdO7P[V_R:UY.)D8f[C1SB,b6UD,8HC=36VU[LAWQ-O8=B2:2Oa.Q2,X+U
[3<2=VL^SfDG7CgY@X[=P(RLK/#(]XZ./C:V75I)@02(3bS>0.L:fZ@-P261YW:=
fde4gF^[>XK\b3.2T+)a\7=#LdAU80FB6e#,A7eIa1S8bQG)=?PQLG.35WYRUV.+
cJ^/SA4^NF;3E/#H.>fVNX4.aYF/J8)-Q-U-T8E6^\6EeFVggDL(QET3g>f5d\37
50NOXS?P74,?W0M1G58@]Yfe;7bQH\L/,T-49)@R5Md3U^f-BF[/^MMS8N&L]A,I
&\5B+7Y9fC6WCRD/bC:^<4GKYOT=_\,Xg_a_JXTcMFO6E_\JBI;?CfGd_P71&M(e
B\-&YU)U1]#WVbV72T=@2dOI1Rd9?^\38RG,H(J4ZFV0K1,V:\TSM?0N>ZegUdQ3
9#[B88&2EHB@[0?3A7:DL>P=WBPHfP=D3-OPWD:[I:)=B]f5ZbE4NPHBV#E^ZG+:
H7(6)9C@O66aQERKcPUUS=Wc.;ON<[+e?KeX/?TUG2.c8287F]M8/MD4NT;NNYeb
>IR74#1&FCW[GN?IcH5#BF-39;UR?Y^P,fbP^7ffN=I>(;U/5+OX#6.)&NOGN:YA
1MW?#RZd1OOIQ\dL#^]N/5T50H9,TR>,X;&b-dK<Sc)gE5Me?N98U7L8V\6&_6:G
)BSOSg,15#-=XNL5<4^^SXOKg(J>BS6]TPD1OLTU/>D1/]-KK@.g]fH2^)RMHEBd
G0T>I641RaEC(;UfJ7U91.dR@W4T1)?I+VDIQ]F._6SHKf-]BAeVTP(336Z[Kb=Z
/(f5K==d\0:->cWW2b]KPRgJ,d,/^Se_3Y/-a4WZKL.#PG3,_A2]G8d8<[;7H68P
_1;Ad0EP7QY+aA@)SXYAbXY7,CA@3(9cQIGe&GMa6^Fe.FJ:UE&d/#Te#3P<@>=L
C:M33Q?@ED+4b/9ZfIS-5#6+;3d:8V[/PCLW_YW@\>1\51AH>Q=X.I:?T),(&S=^
;AUZAQg(HX7<BcM6Mec[>G2246Q9DL[]T=]a<1X&BCN4)D[5Oa^+YJgKMHTZ/9[Y
1RG<_FJ&Y2ORCCPZU:6/W5KN@GEW:#9:V1B#66C,@[OUcBAd&fH<&_KP[O5H60?2
1d9TLE677B&JQKVS78fB6V9N>2@gN;E&I]Q&HNQJYC3/<K4-&dEE_)V,=9>Z?E,V
3LP7A.O(XSDNSbgdaN8?g[EDC_Q?F_Y0DJ3<A1\:AQQ,)<e?F)B4E,K#S^:F1b=E
=&>.X#M?;G@6LZ#4PPd8@DF?NTaCE;@5f9eRdI\57_GFc&.-\GaB82e@Z#?4aQeH
I5/\]JU^J.7WgZ&.:8PaUdg?L8:R:Re1M[>8;\>5Q;YQ>9R9FDMdDcG?&4Y9Q[c=
8J?.PeUN(\NDE_e<9Ug.YJ+1DD>TGd7D-8eF:M7V/I:1XOXS<[ZPDD(W?[X7LTI1
K]ZC#F-@RcL5\D/Y8[P=WEQEbT/Eb@71MJGZRF6,AWfQM3d:I&+Cg#c^D[.(]->:
PDC[+B=<XDX-:0Kd0M9U4S7O\5TQIIQ]cRgJf_IA_&Lc)H_Vd,g=T+MP099C^P7H
ZU?D_1@^+^+6]CCbB-gY-K9S/Vf#GEUP>MYDZ<&(RUf3GV[S7R-Z93OD0U<M=[CG
O>JLDFe.Ac0W(9A188#aEQ@(g=7#XHg0R8WD=^\@,Y+WIg;N@?QH5N>gCQOd3=aE
BASXYa>KQgM(O=#Y&057gLDc(Y;SC8;CZ12M/dMRV,99C3YDca85PN[-aXeZK667
EWJ.&.Ne^=L?:f#\6I2.X3#2NS#K;29-d\3De(&P==)QB#8c()447=VFK@\V@.R_
82NH#;fe@)V;_N]dE9ALR3ISKW]8=?^4I&<I?\]G_gT;OLY&NSC2Y,D2(.TP7T9-
U&AX/TKR+GA\G)e[c)&>,CP@T5Y5e3LN((7Z)a._b=YYKEU4f>d<#0@Zfa9^]X=-
W1EBJFg\_>(cabaIE/dG^S(+9TPDc;ecJC8gdK(9eP(5HT;1,Z]4]deL+_:=31ff
1#32K1:P7aXY5@L;C1[;#b+(R.5&G#K6=d8,f>50@AQc]&#TO&6Q)@&c?b_8]gUK
,<&,.gQ4f;P;.@432UZd/XW^L7=8?H8dQ&[GUcLH?bP9QJVZd<_M:.E8X;I)SA^]
,2JE)DUe<=,57O-@U.XZ9=3^A,RP0@8OUJ@6XWCK:0ZR[+)V53Q+^RdW;:RCJ/Bc
K\-YF<YW_KBR.;VJ@Q]+10R29e2b3V:,4GW=0QOPUCF#RFb\IY[E]f:#,->)_Q5.
W9GPd]3,:&,1]F)XW#KWET3=D&)/baKZY28&@N(^8K9GXc#L.Y1YZ?/O?gP+(>KC
9TZ70,69C]6PK5UP:T_D)?c-@=F=N2Zd)>KV)E3+A-gOgOfb09.4Q</?KG:2Y58b
TGS+<K:BMed+e/P76f)cMC5fE1J8HZW,80gNP6/MD;4Bc/L><_JbDUTD-8ECF3+?
-]),01-:gRN0ccU:6B#P&)YFGPZP6d_G5Q?L7dQ0Q?&OPff2PAFS5Vb4LI#Y]^,0
[C:PIBEOM@TV#-f7)7UG)(SN:-TTN13Y/PdX#AfVH/b]L^WWY8XJY;CJF_7C6)L/
Qd334]<bUWKW4(D0_VXN9.2.-ZRC&2MJfI/JdKRG:OKNT7WAZSC,+E_BST<GcTC5
-P6/?58?e>(aR1YC(bdXM+WdZ59\P]>MMNU+B>[OK]][NV0L_YP1[7SENP+.Zf)a
DFK,C]NGD8F(]BZXC+X6GgU(@99de_cg#XEeWbEJ<eLbR,3g41GZNeNCaM<XPFJA
A:KI-;RA0YaW-;X)FU7TUceOF-^5J/[63&JANb8&]F3dLDcbF4Q8+VB3&4H@cR._
f&GHBNMBF47D(B7DZI:W:M+NTNT4f;@c^3D6=;7)&YS8=4:+:Z,\N1NbJF=XTZ5W
=H8CC&8M5>I+M<ZP@Yb1)5Oc+WQ1+I#YadY>JR>7(c0-4dO40:\Vf3JA,?5eKdQ+
##+2NR,U5Vd?O:Se_FW7/I;==8UCZMWM=&A<NR^URFb_PCA]ePL)>A5&87OD#LWZ
G@Xf3,>6Y.OSYCZZ\FEE;DK@4]OXTa#]U07Jf4:)HDcG&2LN8(bLaL#BQT&-2K]1
IB.?HK53\A/V<(aQ/J<HSQ33DK<f^&.9C4]^0CE1>ZY-2;e3Wad<AGP)?HZ-:B>:
^I3OO#FV+.C,U3J(LF3G^6HZT,<ddg[/?3,XOV>7_b>W@M.]050YWd_H3#W#,(<d
f30279fM,_Pc4)#bT-4D+^A;FW8>Z3,2,<:)J4A&O=4MH3OCe0eWJf@gP.R2&:B_
=#&#3PT_I8;](f;&EbUZ[;B19,P,YggT+I7f,dXR9+>U^V7?&U.87Na_;M(Z,7fd
9R,3g5_fZU#PLVdA]J3XEVYB3QB3N6E8(TYD?EFIEUg@E^IM97<NQ6#VfKOFVecM
(4X]e33Y=5C3^3,X#>cEe>WYba33I/_5.DN,P,_CQ863Ha.K4G:_^8,X>/cO#7-4
UbbcC^=;g70MLA5I]7cQJ^S&RAKG)aT-,:_fD_F[V=8O9;,JS)3?MAF-D1JW[<6Q
/ZR]V#=N9H0MC;gB2O(e5>\@M_YFf,]E::)0OXS0(M_2C.fJGc[[#BK]=W,AY.:d
P.(W<d8^IV6<&G8B_814,BKOa27CaT2Peg^g-P_EQ]F_C.QA]+#2TM=N#a,SW1bN
6e3H8^UH@M5B814+eNEQUE.MO\Lc(L5e0VOe54/EFM/CYB)+OY^NWJbNNTR/((M/
_KaUGEe<T?FN8eb:1IFd9VPM=P/1Sd][^^7B]RRCCKH)J4.^d/8VZ;&16fbDA2@?
?9F>Ece(=QSa_X]IJaM2.3Z=F<SMP+^+>TEJgYW^&<-4:Q4JV]<J@/<KT)DEMA;\
23SIag\41bSIafL=WHd/TJCN)-8Q:-KW]E<IB6MN(^10g1<F3<]WMNA55PM9]g>.
#Q5G(:V&]FF_RE[SfWQ/]K).P@T#,Df6=@(502EX?;KO.-KQ6FMaO=0:Pg?@Mc4d
dc;[)g(0_\3<DIP>(4SCQ]bFbO,6-?gY4NDDee-TS3;8PF5,<^2e7GC-FUaPC)4f
D(QK/&gb34KOfLU(-76Y-^Y6X?Q?5(#\D<2(DHdW>0]H<@3^:>\^D+c#Ba5&gX[O
+\^E^4)A_F)3.JADJX>5bP(O=FT)/6f9f/)OR]E^_7;-fT5<.)[3>5fY02YSbgK9
IdS_40GfI4VQ.579970bR8[[^^3Q>.O^3+W)ZAgVL^1E@)Ze>,(-,BgIgRg>M:);
1?gXZ8C3+Q\<&0eQ7;3fd(_L7[ZW/V--b;Q7JaJOdHGGVafLRUJaG;4/-b^AGfgC
T&-c0JKK^ZO:@FA3(6Y:LN6Pg4dPdbUIP^cT<,>2d0RZ8LScMZ_/X:UJX<I=S\dP
;C_H#(F2)d70,AVc-2^@_800FMBTM.O&#df:.e\7gfc1L\LXCL8WQ6/R.B+b(V0;
J<#c>JXa0S7;QYX.OD&>Y&_S_EcDZ]@(9KPM9_7QfdZbcXcL_#BG91;ZD3WQ+6GS
,@gB]J>E^Nd-20>T(L8UeO,)<,VS,/fG6++PU32gJ=?Eg2_^&>DYb>(STN?-Kc?3
IP0U><,(f1Y_T=[M+#@Xe\IJ\I\\(;I=6)^34Ec9c&PMVO4[J+V,BgO.))\_g[AN
9HP&Y\A-=G]dF(@eR\1JHPY<5\>-D2DJ?>F\9B:1?gZ9DW59aT^DfQ-_4Ag@C4B=
U>M<HSF=a3X\W;_JOe)FYHB5;>daQM&2\<-TW0[@0_<V.?:J<G?(<.@a392FYf5&
623C3<UOcdcFTHT7:X?-JC0;=&?X@L2PA.QdgPGSS8+/V&_-AegZ4SFPV4gD?T#+
6&+REMJ249W2ca8G>J9(@,dV\\61+UMUN0T1&>V6P+YCLZ#Z5^CBWLX13MDQW36N
a4f;Z[9;61.V@HBU(fYDAa33IeSQ.R>A21_N;@Dg^;-X2NY707[c2McCTLU(BCRN
RM)dG_Y7?=gcLFe,M:04&(IDPdFK?B?L-BVcF&X\0F17,&bJE8J=<KQFL/W+U/<E
OOG<HHV)A.7O\dGF==)aJFME#0OTHQ3FS<FG2be^UG(Q>C/@9XH=T1BD&#=/S@c=
ZD,DSUa)UT,U?-X3D]E.DSTG)efNWJLPg2UY^A1)ODGJYI?E4Oc-MJP9M5NKRX\B
:V+[f+bE<6_2.+ZZ5K7.M)2BO>_+PY\V4&IQ7[YI<I[[(Q0-FE&+WC64ZP:H@@+6
0d+IfG0.5H[_.a@KA&-]8^HWTQ?:5aTM6U5]\6E602fIZ;I_W6We@ZKaZYEMe;0V
6W/N.5^Z4&Q;GVgLAaD#FW-T.P3NZ>R2<EP,D,EQCVCY>DECJaI1C9aX-JGe].f(
;8AZ-Ic8RJQCJP?Y[/c0UQMHVY5M.a6/K@?C,95G],V_UV&4I=Z7=+NY11c;?GUc
\6HY,-][e4DRfE\R[3^/N.M@@a#(gGdC>FC4/>-e@dF?a92C^BP:LI4[fZGbP=NY
9WJbE=@fGES+bc;d/-^AAO<2\3UPf:.KF4\?\PM8PJU^g<I/fVU9PF]>-(1@\e>9
?)\>HYUP;OcBKA6,QFefR(RA4?P@+Pea\>PE?&BV[)[H^=C^TA^9O+,(OPBWNIP-
b0L>Ab.V3C-4Q7X8SV6,TFVZ25;0eMOdGgGg7&TFD&?C03K.M(F?J=VISG8c^0e:
(39f_c4,\;/^X@<RCFfT@N?T&cEJN.\Q0E\f:>&/VR_;N10HPWWdHPB,Y-a:0)0#
dR>&0._QaZ.FXTSZ@WT2/0<5Ug(;1SKOB1P;:1SKD1,(M:-H5bJ)C1_U+E^2(^D7
9gE)-R&&.BfaTJFX&RFV0Q->U<E(R?T\01aQW\Q=4X<U=>H6R3-8ID[Z4f#+4d9:
d#C]cJY##5/g2U?I2BKT^UDJ]edK_V_NSE#A&Z,eL>C.BPZGCefO2@_VNV\2PXX\
9CcEERa5.f=gd/?/.A?YL)>KL,WB;g_A74FI4XQ]?JEQ_\Y)D(HcIfCdOFD5fdf9
PZaBWMTeg:Yc<5feYU<<-I^^-LCPAY2O:Y.C48+WVSG&DH7ZT6(g>0),2\RO=^#&
[9IC#4EC&JTfP0a+T&DX3Fe3D&fMg#2a:S]A4U\8E<eTL9G-\J-UJH<C-4-F,9Gd
>)_=F-OAH_W;(9?6)V8(@L-<76TF#D508\A<V?-db+GK879W:#\@W-c4V\#^V4YW
^SFH:8R)VbJ<9Q.;PRKTZ)L,KA1]#.aef.1]+,<MU,@3@F.#.O#/2W)MLLK[9V05
_=M^K[fQP,A&)T,AP,B0IPIfD?72Oa.&2HaF_S9>U7PAVD5B]ND_D.@=QY5KR,61
^23IW)856A[-\gX/8PPHANbBEb_U)T.9cgcTY]R>0I6^PUH;(=4\(+YQ,PS?JQgT
?c+U5.;cUD9d@-S?ODK+cI1_fWb>25O[IV]V0)TY;@DA[Y4PKXL.efPASPXa\@A)
(,NE?U,<&<>=U4Z6O\bA??</b]S)fDd3(O6]+DDBCI>Y5E4HFcFSc7I0[>>-fEX(
U:;Pf#1-d?KX^6fD/E#=O^5S-gDJH>K?,gG._ZdLL[Fc2-Oc+aa567=-BK1CB_e^
LFEO3BU&IR:-M,3FeN:b42\BC?TMRV#Q>]]HD/67X=dC3CS9._38RWUIg]P@G(P#
.+X996e_b0eYEZ\]f0>Q4T+Z#.FB(T7.)(gG[+XBCJ,YZLH17-(].L+IPF:dRgNJ
T>O:)#VL&CGP)9[V(XH;>f]/I&+AI):N7W_c9B+JX/X83))]HBYeS,&&I)gaB5b^
Dd@YD+9WC+<HMP;G_:ZS82D7NRA2>5<=2<;0bL-QQY][>[]BL[80FgE,F:0:?3[)
=eSCSY:ZJb&9+,/WG7\:Fc+ZJCdG^53;URJYEFa<Y05<5e1,#aK@^&^_Adc5BR(X
DLW\>NI6S+BaffW?GY<X=8@>b-C8Vg8\^9XT/SRD,1g:;0I^/6)&ZH_ONc/7aX@I
;#&[EQ<@9;33?8V+]743JUTg4E-B<2\8H(A/ec)TN_Z7NG.2<RaO,)cdH?HMQ]b#
TTd\\A.X7O2UU(J+#J<YV;6P,M^W_9SYJ+6NN7HJ8Q.NQbd&Q/_\V5+J-,;IgE<F
2H2WRP2f=,H00QHC7(\:KD0fL+2SQMT=URd8UKV5W)30d6B72[Zb\Q:6LX.J:1U1
e?S+E_)P>UD)&Ka?Bf5A&?L8[KI[[eWXE2#4W)G=7;J&gT2c?^(NVgf.B^4_X^80
2L,CIP[7Y2[FM1];PXM])D;U5&ff.YALKEgb:<1UF8NKFW8=JY4J.C,_XgdV1FM6
+F-HX>M7]XL.0G):6DN.1Se<K#0#1[@/5L8KF?^2c-8E&PMa\,CA]:BCW=gTa_gH
^O7\&bQAK(:Vf5ZCQcaUXYLY>c48J_.[f(eAUc;TMC-&57\XGB:-H?@D2W6B1eQV
.XB)a<b2aA)=EI[XI-8>A_3^V5VZd,]\40#4H)=g:afUbT>V4g?08CE6.N=8@MH4
G0O1XL?Ab1=CNWa(YELYN5DH1gU^W(1(Q^TX,.5e=1bf(@Y7M:SX?DP#JPIbCRNN
,2ST>e,G2>g#LB-cY>];NXKaRPYUb&P4c+68RWT;I?baJcgAO(>6R+CPZd.^CXH8
[cE[)CF=_MV#(&8R15LK,g/-L[PLa>cGX,a69PI4Cc-1+Ee(TCALMUS(\<+cc;?)
]4GMeXPIEY18P0NCCSU#<&gU#KHS/[Z(DSLZQf-R-K2W2<A3\2:Y3_b_HEf_3:;e
_Yf&/[0]N&A<H\(eg7[QU;?HKI\..GHBGcHLCg9JXa:RE0ZY)R09=0]H:\DCQG:[
Pe5926M,]5=#6SRgag3GZa<=\:KIfHIAfFD5LH>FL7-8WS,I[42EaF)JOa#N4dR]
K5.WY8#ZTd5f#&K&e-,.F2P;L&8?W/T#aN698>9fSOZ\d7a6\R<:WWc,@5RASHEZ
PdLD_QaR.0V,FTF9[2aST+4GSaM2L=IG_Vf<:;UT-C.d6_&/g2NC6\AT:=aV0J7N
4.=)NARXODVPb6UNUDMaC)3]BF2,M1HA&F<d0M^#8Jg;6cYeO2Q:0L8I>[:9^LL(
8,EbdE^HANGVN^d@VaF\#2.45dg9-26b0(SW:XLQ@F=GS/L<6LF@8ZJD3eZ;0Mc;
C6^:EG?^:f4::B(0@geNZ5V[]9I&EcP0<]\K&U5Y&U?G0O/DA;2B^\T7FTHK6C\K
NV@_b9?\3R9:E#P>[Y)H:a2K_QdX4FdA0JF,g^I5dG8GB5+-#c0WHULWJ]4SU^]B
&44./Rc=;Obfd4K2;/]T:ePHg=78[ML^S,DY\FYY]?[d@VGQD?aYH;9@AePbYGD.
(W43,=63Q>Q<?4.RPSc?>KWRVQO8c-D(F8F@LO[E+g3AEH9)P2OO-B6CBP,JG:WX
FOC?\7)FC(A<OJ^FcTORcO0PL[2E8SAXAW<Q2a:FGY_]a<Z^#P9W5IGHf>E@4PA,
1bNHeRHROD&MJ0CaFC.f7VRMNO5)N1KP-RO44O<FX(-Z=0e(TPE+Wc/9<]X2c[8b
;J1MQN<SI8?8Da(T)@J]d:+UX.T?(8a,8YR?.V?G05O=GeNJ#<4YgR-P+PLDU8J]
N,@g1/IACd7bc<ZTP^XWIW2(TY]:@_S4b?+GbCFUdN.IG?U<f<D,:]8aO[L-e?SP
\Bfb)G,D2O>#7U9;U.-F0Og/N/bd(VPITCd3cBf(NV4QET\;G283+E]Vf2QB2^E_
d]UC:+Ef\EBCO<e&?e;Y6Kd9S84<].ZZ4QK^-X,IGI?+1[b_42J<Ld16?ADU27O^
UIcaSD2-cIW;O8IL(9_9&MEe>a4X@3J+#(92V@Z:&g3M8a.e:c.3JS>D/-M59g6X
@+ED.DZPA7BR5N+RCM:,MXR;[HIKd&3<b6P:5,FYQUD_PgZA4Za^N9+:GfP]SX/M
K2&^O1ZJccT(YQ(.5O>^[TJ^_?;(&R#.28[C_2bAW&4VQa7@@L86JC/6>1JK^2(R
1f#,&(b@(]-(_WAaPO?fbO0/b[DK4E82g2,HU>&(HfdB/FS2],gT7:C_&([6L5c6
RFc59PD#8cLAAA0A@>dd_K8V)EXBM<(N1]P0PG[?[Ja^8Mbe9\P4b(0+ge=I-0N@
.8D3/<:Og@G4FcI_[1JQ@B/Ib[Fe+5YZD^WOE_,YX<=,bY4<gC58B?9-^R/&3?]3
>fc:6H-U&[&(8U0;)W@(ffNSB3b2G0R=&g_<^:fEMBA:@O1ZM,\e9#7f(=?33^9/
\?gU5#BA]a3H(WPSaU=HT9#B_AIEbTa^1#Oa06Z?IQ#.f/F9O3O,KJ.U<>g,_TBX
O62&P4>T4\7>CPZ\?J66@YM>e^#\g:CSXG1:6:83&31MZW7X>>(daQY&fC;HJ=d#
+MZeEIeYaf4+0C/:<?V>NL/@>T;>fPLZ;G)#]Y)VKV]RGd#bMYgC:-K[2[NCG.L1
V+9]<8\d9W?[H/aJcKZO+9-IJQ,R-;+#ae&025c#gP0O?Z)6WSRUK9=/a31)BI?7
T>Fb+)M1+W/QSY^F5S]bWQIOZ-<g(Qd3L@93:+^g^A[A2Z)Qg\a._=cJ3P,eYe(L
EBg>Rc.J(=I\XW:^PQf16Id+>T&;_[a)VR3_SGEfCZ;[,-8d]T8@)CY8QG4+;],/
R^dg/MOKQafSQM[KM3fP31Q7W6AdcbS+?=S<V=JD>-A_3+a64U]Y=3_XL=8=X+KK
N2)UWZ:/R+P1/-RG:>\77MY0J^1VFH080A1Y0F#6Hb__RSHZgK(S)(a6C/NeaC]S
a\>d31NY2+OW3,9F:Q9C>D_bXKR>B@7T6WEe;>MCLPEN5MVK-GG9L>bD>;AY)PdM
A)S8,MV.#>0+<_-0ASF)c]\Y.&I&CJE3PJ=4SAH^C6#QS:SISc(:VI/N;XW7]W3C
/?e:V\34^YOPMG4A+:EI8I9IEa?)KVTQbKQ60+X([cQ1YdKB,6_f+.@]cCGe,1Q?
f/\N.a6g9(_;N2NcO5^6DOQfU3FZD#R;\)=M4TGg&bNE1d[-LY4Pc1\8QE:<-=OF
0ZLR:Ge>E,]JaWV(5I3GbCC@;KP/@(=4\=00A27Ie,/F-\,D@_;X2):fJe=Y9(eN
[0fRPL6GFKGBG]K2(I&IYf\QF9_gCQS=@4eVHab4J#]/NfaaCgZF:L-QN1M)C:aQ
3Ce2(FZ\JN41cF9WN<]@<_dYIf==cH&3-\OG5fF<A#F^H:_48aQSR81&/+H?F[N0
0<AWfVb1.E#^WYS0b7[I[Z#4H.BBFXC6=#9JcV?YHC4Z_+MU][Q;RLDcBT[0UK1]
AQg0W^I0#+9_WNeW-@Rg-aV93:JN+.MD8&L8</O.ID]d/Q[GMc4DCP^?XZD4S]gF
geQD79/d,]g53HH^,+=T0_Xb&BI8,5U#XSgYQa(I9M,=@6K[.&,1P+([VL+<A;K#
^\PPG>N7VYDX&7gC/>\d,EM2&N#=8;GF#[#C@UZUGHJC\QF[:#PQ1Z@Wg>,GD<^9
2M8G)M=&0DO7=b<eUUTI1KeT(P^g:I&-ZBWMMSfP9@3;6JBdQ]SI8dERLdI5g0+3
JdO1FTV;e2&DG6cT28-.FL[:YY6,T#;eT99H-g)@Wa9+XM:T<:W\)L_cDR3/A\K2
^g>X@]MJ^#<8N2P&(OAOQDRAAf>53)TS[B26/+eBX2X#.GV0d(eL[A>5Y]+Oa]U4
DESL@,R?_e[(^G]+U>PY2&F;R8B.XAePA:e\@d[7?P(EHT),[Q+^-d//ba4^(+67
fZ+^4?f#G):gF,Bd6DcK0Q&L0S(VB36A/C)L7(6XdOQg9KN<e<cZ?/5K&NGV=W4V
O92)bfJZKCYA7=KM?LWJHYVSQR2E=?f>[=DJbXNK#@>&VNXN^)/>cf1<DYe/;KR@
IZOKQF6@/Q7L&/S8a[\IRg98MV[,8D+b<N_>e<^(IXdJ@QD0;UYbNc/V/2[(P\Nf
0;-0.[=M07-]&//Y+D7=E@VS(E4>TP<1bJX:fA0\Y0-X/=cQOF<_,BJgbPaWJdb4
V^d9=E;:UdK@5/YJ-SfX\FYQd86Z]Y4B&5NW.1Cg1_O2T#b5MZCI)\[^V4Oa)ABS
)1S];?4INK6Qf?]L9c5VBScd3_C.E=F1P-0KUI\C;4/P7YV_@]V=O/&SY:aT9aI1
:9fCHNEBIRCWQ36Gg@9Da=L->F(VG]e.12@a?[Ob@OAUg);=]#Z7M10-Se8PEC3F
I?64QeU:&LK^.8-dQPJ:.UO0Ve.JRX)BY8/J3Zd-e;:FB8AE^:#&+WUCPUZa;9>.
DO);#XedLIM>f7G3L8IO:acBGZE^a?U^\P-c5C<=:]_N_KG[P)&LLKF>^ZJb26__
4,PV\g(QTI5RgEeYRZb+c[QLEbd,g?=,ZV@6g-gO#GA1\=ZAFUJ>\DWB@]@XP,Q(
_77d0,YY?G[S;OK<OU+8#:0?]fWEJ?VS?N,HH2SR3LLQ9f:FOK:8f#60?BWSAFH^
85Q?/JI:&@T24+TG-acb?R/>C&/BQe,SO3[E8Xa3F9.]fUcYPM2TP3R]5\JG&c;<
@2B3:BM99Z2-HQ0I]M6U-2bG@FeWbQgU1\=OgQ(G8#[c,MINMW6EI\#5S&c@#Wc\
J6-HN\G-F5g3-D9(&[ANZ(0R40GeZK0gbf:B4CT@V<\1QUD[FD@J[OEH[W2gD(B@
a4E/:&be>-HSM]^_:2JXf)OEGA3#&>PX+gY+bUOCUE8aCHL6XR+g-5acg/;g0&9S
:XYPK/:]530NRGVTbDFdQ>=[dfXZ3LZF83fB@#0M,GN:JC84H7EROg8K:W076[U8
86:Q7SEM.Z]IB2X2Z659K;bXY]V]>7DI8IFDJ62;76(85EKcUG+&^<R_CD[][VSP
&M<8+SW/2^fOOPdQ5F37#XdY&.VK8C>JZ>#T@KXS_HN]::S:J;<PQL@N<MA@B#UV
,<?eYZ0@D4:@ZEIO:\Z1<KV\/AFVAD#]@E>g4g7c9)&,22;C:/<_;E.7:eSOEQ\M
=W8GLcL;[b4E?8?1ETLa-I#d59EB,F8]aJRWGIa)W;R7Pf_^H#4W&2)O<\#8K6_>
)G<O6+WGZ3f+6Z1:LR1#+KL04?:986K>a2-;6Y.BB,U/D+,8[b5X59CH48#SAdVL
9YG3>7VB:_D0YHeJ-0\VR?&H(-eL^?<3:(edAXJCe:ZH/QYbfBN#6T34c:NBKI69
=WIF>IH,INM,2?)LO+e6PRF(Q2J0I[+T<?MFR<\dPT_,HFYYb)/BQ]H0aNY@VU-J
^2Z>(D+.+T-_@PT)bKLfAZVb2cY/,RT1CP\CGU47]Vg>FP7VN5RST=XEd#LJ^c-^
?4Y4^H+:R&X:]S,^^-:M55^e?MTH.RJ42f;e@)Q.7^Y-:I/:#_,&M\d[+^-dR]RZ
c3?YA]3UHAXD@8e7VO7(.aBUO]f-1If1?W8TY18=aU2SU2P+D^fTF7:U-C8U<25T
7J+d,=VLI&HICec&4U6a4faaegHL4ZQFD_SKePe(+dCA.IQTL-^NgO8XS?\ZH>U4
eUE_>#QS(M?ac?3+JWBD0RfZe@FWeg]W/:H[RFW,>ICC>6PIWbR5ebF@[K1FX<77
UT@L0:JeH&baNTBIL1cGA=2e&A_GC[b3/Hb1YLGaZS8[d<g2B99[:SKOfU)6YRa>
CB0e,<,,/Z]HCf\c5I#+LQ8V&eJAX&5:3/G@;I#:97I.g+WD:4#QSCa81YO#8;Z0
D7Q.;f/QHX-18&@SJKAH/#(eRQ_X(1;G;fKg2)GMZSO:/D++g[^=##JYL+ZXR&G:
D7W6DA1<4]d\?f@[V9La]LGgQ8geMeEN]N6f0NWSD56d0MZW-K[5GYb\)\d[(D;E
Z<N;)KM)?KY3O4Pc;_6UW#PSebQYb_a8FV0EZa/g+5,Ube&gLg[2gP:9T]=7gXH7
aJZ47P#34TR;]3FTe2]?e[e)bKEe9]4H:K?_HDF,TF(4e:^4NVN;72c<bPPJ&^a;
e8,WHB>N,R9A5Z&0V?OXAV@,8FCDdLOYVM)__^:HEfQMdA^_N@4bF46<?HH8M.^;
N1Y;H423cFFV8BE9-K,W;W]OLAg6NK0<)KKZEM@/,QN)9OF&0G2XAWQNRbR5>Rd_
\bWZ7G<J:\YT:Z>[WcbG7MU8Y8LE\^78S4)L+<A4GG:@,(U/[W7&N+LR^/ZMET3+
K+#1KdC[C^aBID8f2K<]_1]=[S13.\:2<?WRKI5:&H7D3fNN.4(C.&9>SJ\8Hb/c
_Z])C5c8cRU+9;eQPB#Oc&0/VCI;gebS?3-:JF;\TW.ML[?J#?IJ>4O6I=;=_047
[#+7g-.ED_fWUX/RZ9O3M<;]45IO@@BL]MQXdG[S;OcD##<[L&.M9cNGY\3C?V;A
9I)4A-(S#D1:QO2#QAE_&&+Ta(-GUc:AE)ab^[EBVWAKZ8ET6+@fPFQHD_35XL])
RM4[(\gG4V[E1-1@CD_0#[1FC=2(W-0EG37@7SG_^VFZW:5>-TYLH?EDK69_b)/0
YM53C+fC6XJZTOXQ3?E-dUL9#ANY@LNO_a@M+8A8OX^.LG;D=OUUYR]E24X>[Te.
F5MCdL4\UI+bSeE:IRK8ALL(/#0-^g-2:52J5>EUD=130H^IJ.Q#+]B2T>9FSOPS
#)5;E&\/N?VUca1\R8?\L_Eb#8E[^]^NZM-5=W1]:<6a-S2],>DX@VE-5ZIXAc\,
)WMK,RU6/V&f[UR3Jf((eSDK1).GFQK&=)#7C0(;\U9Ig,^6I^GS:XK[/LbP93V,
LDLA;/?)DF@a4?(/DCB)>e]/)A\/LOCH?[B:16:,6HK,/S/X&+JF@R&JY0D79+4X
f.PBJY@J-IDP1KDGf?X@R+O#&=B1A[4U8N+@C/.c2/5PI,\MZ^H>=ZJQ<2DKWa-B
3/YQ0:P1d4\2S>/.<N#((9-:.LeeMgH^LYgMM^(^6:./S2K_^d)OP1P1dac@bOGP
=+-ga-Z8BI)+G&bIRd8(E[b<J1+dgL-18(:=?#b^2\-Y.K2>E8>bP3.H9(;V-(fc
-_=NLJO]O(a?bgFSICN2PLS=a,IL^:[T=+:B]ROA?L^Z8-O?#_e-;YLbA##dHHaB
/8NXX<_,J-?9Zc_PUECg:G=3AUNNA7NQ(S0S;_bd@dR7@]UY^MNe_@U4&M7?fGBe
TT]fIa/),6+@=HQ^:;Z5X2<3I_8C,;>^;=e)B3FX>WVAb60:9GOA[):e,R^Y7\YH
?/G^\;f9Ce&#;/5XW4G-Z@F,2a56QEc9^&J^A[D=O6(E]ARf]e2B><a&?UeO[Q,W
f))RAWbNf2P>B-]_)a80b+Lb##>Jc[[</]11&IZbeSXYRO([8?c@+.@NC,c61S^H
,PP@92\0U4PXc^T^ABdRK]L<>9L_C:\,N9eZd-KHUEED#e<[,[)3&97E5HBgPeLE
Y@W(aM7\#SH\G02e.<6F7YgNeEI;?;([C9<f3JUX@c7:8\M_E[]=>Z0BA8A\E,3?
&eWREA:R_9BLC:?0aI>-=+Red15eBMRMT_IbB^PI6ULcC:a-@971IKF?5-f?QG.W
GB4-]JRP#IZV[57EK+G_58?DfF.Q[;d<2L:YC7g-\T,YTLDN[:If^6fD9Z(Z2Rf<
La&cc_1\BGU+9/0.[KLLg.fd,D=UB8U0M4OW;LUD_D,Ted6;bS_1>4&Q\>ag_1-:
\Q_3,#4WSI&dGYUcM[1Yf^;_Q?)K;)9[_ZeebS=7dGM#&I;.ON,:W33:=O]ET#FU
H0O?WGXd19f,#=_e#&ZKNXZ#=VN5d8)8F0BYTE\QIF/IDdJ/d@OJLQe0954_PCbV
6<D4_V60:bKC@a_R3].L[KHHVaX:;05R+)3#H:O.=AB-XAZ@=5;V4XN2_Hc5-:XH
NYZ.1b;4SELa2NQH)RPS;de.9L1_4D3((XXB0+eZbGG.1^A&I(b^F+887WX\Z]c8
8OIUPUR.(f2_BS5RG1g^b\J[@U7I^E.#ZB+45#4b14IgNCeH_I,=ODY6;(SX;/OM
eEf@Y\LP8?<C?SJR1BXEK6IR@IYGN+&;R=B8@/J<<DB4A+O]C9d-2\\HRWUR8O\0
X+@M-VP?#&120X;:.O>,67\P9@&3.a9C\]NV\RWG=S_PUe#N+GYL1//^6(;PYPPV
L1.9bBA6QbddNdO5F)3Uc0BA2T+=9RS-S^3T((9R0]8.)?19E>M3:Qe#L?cXX3GB
V.1,GJ\Q)OLZ6K;3_YG(E88fX/MHZc(5b.Gb8BUCMQ^UO8WC]4#+>X^E_#034K_0
E0Q(Rb:8I>ITYMV,PHd>IE&>5]V\<1=UGVY5T230ZIc2;eAR;L3(SA,,C2@B0]XE
R02MA^P3SeJYPC=SdP5\0\:;R19:,MaBAWgIUFVK>QOLBEE_J.Q[)511C9;]VaB8
+_3aE[-e)T\6gAKb3BH0\4#/.+U3;CM&33J4[,BHfd:AN5VHegGCOO)<COW<NZOC
2c\]1YLd^KdY31dgK?1>aeH1)MDNeK-C;6AT(a)P14:^2.+g&?Kd@ZBfM^FAN?=B
(f:ZO-@3:DDH[,+:N7AXB/(_=8/SXWSVJL(,X/5<PADfNNNgUDRQO#Q;+(Ha5Z\e
.b8GII;EB#Bde@Y-:WfLE]_Y6Z_f#<&],\G2T[3CZ#YZ7HXK7L4LT],CKXdDUL[]
?]S.,C9d]KJVV_O>^Uf<88B6LXT\aNOLY2aC[A)BZP8;J?eXa9_PGM8[g^XG8Se#
=DZ_=9N5-R)<WTZTYEYN<]P:]&deL323JP8#J/WNbRPZRg/4Xe@f:Oc=:WO1WFH2
LC(KD##V&>eAbB8I=BI1#6EZ3fUILJ>\<Vd;S:Q7d/=)),UB/XcFHB_f&E53NKDF
VSVa3T)d]/J-O1ffa>+Ib7]eEVE_QCQ73G)#NcBD^c#IdS,91@Bea3Hef]5\]AQ0
P>PNYg_90;9FI3>e=M;;]+U].#4X:c>e+WNXD:FA#IYccW#0GBS3>4I,5M@a6NJP
K?XA[>3C_>03c=Fe>.EQ;0XOb2e?;K\0Pg@0;(Q.Z<>.CK@45a\9:&.2/]-.RXJ^
P6b5T]F-d/GG]9)AHL#6V,gN\</ZM5HTF?c_8TB9bXdSVR_Q2Z(0::T+P08]?TDc
>1S;R6Ka#HdF2ACG3QSbfGH],?c_MHeQg,+QVS9UgXJ,(BDHECVN=U8dKXTLC8V:
:E&STT95Z<I>3LggLaV0:<SYR@PT2E^0eA-MK0#ZWB?#T09;@U<0H8de8Z5\ff3E
60e+F4IBNRSd<+)@X>58?YM[fA4(UJS(HO.=]+d>>e//?/X/MQD68c/_;B9c4gUC
g3Be?Z/>H)0;\QHgJV9WFMb_VRD#^M0WHTK8@+8JD8MK=H]#.X0^XcS4E:f0H])7
.bZeMB>.\IH+H5-K?aU384&cV2-e?Mb1&=:PQTAO3O4&R,;B2)UVK^Y[^=HM@MdX
H.P?LHZOVSUReWL,e[(3Iae?BXdNbf8P>;S+TbYO0^,E3:O<N_C92U?c5WfT>g@+
^e(NA]AM_f7c_F1#U0Z5VTb5ecg_7K-;OAOG0N3215Zb8S5ccB&HRN^a75TF\LY8
]\f:M?/JUD#3RL<g2_Qg+416QJ2cIFI->T86g&)7b02D(=[-:E@8/]cB;ZW\/0S#
M;a=L+M_?#b1L/K#2B_?:4B(F5,f)>]H9X+@<^Q(JAgJ]/?7HD3.g.LE<DPfMgVL
NNJGUUgcaHI9A_RId?E;T5]9?@/K]+<[L]C_:Z+>\UfU>Sc.]O?:Vb1a2;@[\DN6
:T+U6\EVS7D1&PT;_g9+NW1Fg+7(VcZTXU))#=dW.EL-?g@f:VXJ]]:[;^U2FTdU
V#+dMVF3=b[R,-,D])315DPadVV3<cZWMIdF3889UX8RY?F2;\S9>)7MaWM6^?):
-2#8GK2RND=eBUUHDG[D6?8;-+4a,:QJ?a[e-TAJ/DKRYPL1QBU,e>C]8D>Xa0K?
S//(<QZ8&@KZ,ENLZe,(C#-8+O6=_&BS7Fc\/Z:MV].6N5U1Q]&,K+==&0J)GG<&
,V<5\6LX[I>2YHfbYf^X_5N](eB8;8^fQ-^R;?LFf\PZ24S=0S_,(bQ[[>K(6[6J
>N=]+;FAVR,BDAg03C66Ib;@=<?06N0(2CW]ATEXMIYa1TJJTCGfAH#2K1N:=W(_
2WC_L7RKC42dWS=7I[\<Q&/bX?;cX,46;c9cffP^F@I2JCZ@T2L9UGDeN+.?f5RV
J/GYg)<RMA96(bJHNLJ-O:YQZ1]2YPWd+NX8,KHY4d@d>#7EHeX739B.aUYOAa5_
E>b^b@[2NUe?f4M^3;a_9ZfENBNWVSC[.4YDA_<B&#DBFgRd&P:\O_#C6AJ^N:51
YP8P^4/EO/W=PF^R=A\_4)3F?>SJ+@LU6d)]gXI[(+R>XV?gd]:[P#,f99eLa5GF
:PATP\cG+0EFZ3^\Zga(QR;3N@H(877E(bPR[;gH4g<4IP5Q:8ICH#2H#YcEWfKa
,IHd(Pc7R/3fYGM9_G<eV1HAQHQX[gQY^Y66\X(0NU]ZQPUNKEU_Q;3QBL6V5JE\
S>W.-^?::S#RKeS>GE4/bNcH(6_W@YKM1=]^,/b+I3GN4PG41&XbKGJYeINR/U7V
Bf.Zb;.V)eF\?O]Vd(H\4NGQ55=U]EV:(JU+;Q,bHKee\(WQaD^Q4F?GM2G)V7/L
>R@I7L./&]5?NYW^a<F@;(Va-SNHPGJK[3])W+?J?P@6,65F1YY>bWeF<d3+8W/,
cK)F?FXDXG.?ZK-3),:^1gJ(?[#;DGFN76JZdC:FR&Z88;T;EQVO^VRO@/e-8?g>
:(I,0)4[&P^.B.LBf[-J@ZYO_d#cZ,MZ?OQ^M2PIX(4JeK304F_PCREUJ6VMN^_6
7OXXBL\<])7fYI#CT.;LTd4RK;B5EZOX[]Y[1],-H6//]DP#e+Z.,73WT(0I0TRZ
fb^&.C/4I,=B&XLgC<ZMBH2MbAVSQE=>1P4D0#fMU6/2<]OB@fPgXd_d(J4<LD/d
6Y.1GWI3/EFXg#B&/Z<(&DfdU\N4_55CWYQS0K/0Q2?[aAG6IQ-.;3fcF/_Gc?gE
UNP6^UdS^dF>B<L);Z+0SH>)T+#Ag0\SeSKF-6#[b..<[FU&gZ5f-X-Y<>LgX6WY
@aOV?,UY+UG+/da:;f@P#>4;^6>d^JX3EQ9=e\.8eGa#aZQ8,d?>c@_KEOgXZW.7
+W7.C4URKegYg<4cE1S_.CM)F<HRG7S=X?g6)b55Uaa<45\Z9(KJX6.7F=_9@QC3
VH=VKg9GR>3ND1Td^ecba&?Wfe^NdA:4S;Y286HF,CAUEQ(K17W.fMMYX_4g9-ST
JK)<EH=KS5WM#aO:1cOWM690+cC;0D->?MZLP^G_=DR_ZMGK2HWB_+8B+:+U7>5Q
#:J5^PM2I_,UMf=KE;eVNeJJNKeR]5.OE=,<53XDe5DDFeHPF_9M&WaLF^Qa]8K#
M5=ggPI>5M[4cgaPK>C)g;9VB>1GgJ#EO)WVb.T\a9;OG<;\#Qd5Y4LdD6)D5S/E
&_KR^c5&^6V0cU3_]+N7[AOY=KEJB3@DXS^+Q\3:fS>]f?8<U]\?I,SgDa0XD)Aa
Tc_NAb\b0_3)#1AC(6T(b.5\/,T7.12QC,e;BZ-Xf::>3#]f#D)Q2U5X=-BYgC2T
W3aGf6,78TO7b]JT)),;#[#:[_J45=YE=;/9QgbG;POQ_J4,VV=X2H;)TAKXCLQb
+[4^>,-DCgBC[FNYa[AbJ]B,7D4+YD;&H@&dL<A^:Nb_UEIdI23N;BQ@D,WKac?R
e81+[Bd]5MK;b=Qc)YR=IK;D>YOORBRW,=#gX3F3^OK^&c<&8++ON2Bf^;RATN&X
g)fKA+N_O<dG\N[#3W6+Ae[6KN#SW@P=g<SQHY/1UeC-IKOOGYe+gFX,bJZLU?Uf
d/JAT64T>5_+bP&B[SQ1dg=ZL:)XK#V:fS&Z&-#.<aMbPeD?G0@(T?@IR_QLVK?M
[ZfH5KDE/\bG9D=A2BET)./aKVQCGN84<\e;8_9FS(dFYDH;+<^CDZ&aZ;Ne^Xd4
[HUO>9[&G6Q\.Z0]gQ0McH:\.(WXK-SR[6MY6,#I[N()T]3SCe_PJ?RM^]Yf18XL
1,F2=,X;4C[)XG8-.a_.\MKNIS\Te9F&2+KN_;H;YM:GK:LQOdf8V]UYD?X3fCd)
]b+)=B#[ZL+WZW6BM7DKWB:,Z\V#TIMTcX<BGFZfN.\7F]:dXeWK@O-b\<S/1&F[
#dW@O7AeT;aDGDd\LVX-K3>7)-(C0CdJ_2DBNf(.XN56(Ze2MDP)[0=-SDDW7^HH
>6gBL6_@RRSD(;F2JKXYM1O-(#V?-WK#[NZ&,5?)#b=Wa<POT3GcCYSX-g5QdYfQ
;]6MZ3P)f@[EEeAeMJ=@N8+:.R;OG<.NZ+7J>VY.(Y2dd@Sd9ac^300\4,JUgf@K
+e>g)?a0;A&R\3AYgNMR?7?,eP5DTe-4MJdZWR/B3PYaJ#\BcM_DE9+EEf[e<>-6
gJ0eWBDF]A4.f7eX4dVQFY#@C,F;FbQM]H9YBVQ6GaX054><P\,-c\QNCI[I+[Gf
TX#a/K-I4H)UWIa=V1Q48[9E2M<V4,gLgNFcOW7a98Z9:\I5LXFdGP2AP;BMVS50
e&Qd\g5U=^;:D0.0+U(ZMQY,2@H>8I4VCHaOb7W_HV(BQ,Z);QAOg?:Ke)[6aKDA
PPO[[//&#11;#Z2))2E)DIXBQ75<RWL@ROR59AD]XA5,)@402X\OEdGPRKWL.c^@
.HE@QQCH4&]8#R.LWCC4Nf5S],9VaQ&UCg3edVLfAN+ZBDWZ.5[(V)<GRBSLE4:@
Y1NMRT0@OH;V51A[N(@2AGO=TV6.Pf&YG21?=?Q&ag?cF^8C)^GJ[FIK8P(6.74R
cOU)FAg6?PSYG8Ha0OTI(a[Oe9K?S6<faLQM(8aF.5)b9J(KDJ6G8.94dUaa1\D<
PUQJ&SYD..\B15U&>;XSI3c]1&dIH\&2VQ)2_bF#9,Od8IdB@^,.\d@E]D;-6>f[
]ZEYG^DLB.C;N(B^(W&VP)PC]]^<U<>7THAIXM@30WQP?M.g+R3#JX2]/1:fZ,(\
2#J5:ge4NOT\]3@56;X_0<dfWIO<VdUUa]51W](J]_FFKd9e3[_SUb@2_-1cQ+YO
YS^(cHOYVBK.KH?)N+ZI#N8YeAecaGW=R+4.8>#D4B8eTD8]?U-;>YH6?LN2</6?
(MTXRgX3.+=1A(VHc(F14)N?\HgVNO#=W9L\[:f2dN78<FWT<+X6)+F;@S:aYKMd
,(4Fg2eFb/SAHa-FO3g;&e_9=GOSV#>P/gXM+5Z\JMGH^&)?JM6d6>L8ce>cW@CR
-eXMbJN.&Z\UM]_CCY.UXHI0<J8L]MHF&^1N,e59XGA-]#dAV8)K49MPFHJf,_W(
J^:-F<T(9gB@0,P_[94Y+SIGLPeJc\DaH\Vf^+GIF,[YE#7Z82VES-^9cHU.X<H[
+T;RB(7dRd>XQ=\P\R9?DI,@/<IDX(OTCd5e/Y^gR5R5(_G,9SF/Y,=\FCI(P?,4
Q?O<^^WJ:SJJ#UTZ3Vfb&c\](B0(6VG?>ZQDVEY[6=#=9=>-10OZAR0&]BC+Ie<3
>YBW>.;ESJX):e1I]/QH>P12#dWdf(WPK,]2b=XXfc<T<1=+&38=NON43T&?1[\,
Bd4I=+Q86;6L#Z&4<]3N3-FMXN^Y4O5&cffTZY5b_PgcX2>d:XNP(L@RE_3fE7aE
(-1;fQDg7eYTY5?B31\SRK;JNYdd3/D-CQ:)XBS2AP&7)G2g)UC/YaGPV^O1IAFZ
PVTZF_BNWZUUZL^JQNKZ?X&YVQ.6_I5MZD)+8F+.W<TDN64g)g/0I>1_:U3;JMQg
0db;?A+RN4,(3E=?HPAF,.J^PY7?bHd7:-Hg=PV?S\5+Ng3De9.RMLN_&F^X&,c&
eXXfFcbJ._)JB.RTVO<c29&6_PYEf=.dd9;I0LRSf6B\T](AQ=(d0<:M?P[LJP4+
@&@?K(^],\_0X2/UO/X[.Jfcf<TNHWWW.Fg_gS/C:R[?Ia1fWK2.EG=d7M[J;fGH
9DM\M,887]:c&SHbY/Z3?K6V9VANcd9I(BJb@32JC9SL<AD3D9B)9@2E@9@fY;c/
Z2&eNE5fZ.R<S(gag>EF.-L\S17P4V,d7C(S^R3V@W=>D8aT2UaS?[3PA[6(M[\9
8.X4O2/=Rd1]I@X7I(BH\dTb-E9J_\;NCI/]R18ZTPI4B-_<d(-JcA4d0EY@DGK5
74[AD^dQ/KB?J,&(IO_6dPc^6,X((V?c^[D8=Xa_c2+]?7deWYOf>Y2Y[9=F33c-
;&[CbeJgY2,VCaaSJX1eZHL<PS1)IUZA]J,KO5OJ/@WQ?1</Y-b00>:W3FeUQf3R
CP<HbC;OfYHUKM0K]XMCIUcJ75JbCHOY9I&<..3_?<61+-W3T7#6?LY]R#GaX[XS
:4Aa&),>B[V5ab0Y[3cXS-03<,@9D,H\<MGRWNXDO7c8IUMIXT4B+A;M7f0FF7cJ
b+<I84(LJQ0ZKPF[:X7eD8eQ1])58\^>LT>N;H._T/XU@JBZ+f(8M[E=)@TW(R=9
=EBYY#-F.>6>DXG_VYZ9KI-?5IB#T#3Z)E_dRFe0-CA99YCT=G4A0a3P5DX-Hg&]
Y(8f0QBOW#c&U]/J#C>4>AM0Q;)Ya-6+#L3:RI)Ef9H#M@N[90-\XJ)H<0TW[B(/
.(?,(U\8-]@JFC2BOWKRQ#[J63:fPSdUP]L?_-B+Za(&[b>gb4-Z7R7\AWc].&dT
2(/2N8CP#5Q<;RPVXSRF-W0XM?-ZN:M<31,Z<d?[I/<]UX@>(fGA]8]=,=g7d]0Y
B9H=0X)LGWaK.E/R[JFEN/MUX-LQ@(^GU^4;-EC:OFN:@:D1cgU0QV2DI<9Z,8cb
a.4Q,H:_()_=:--8:6:eC\X?UDY(6S@GIgeSY+SG/=7;ZgTd=(;XVU:7ZKW28K5:
LX=R?.QM17Ud[^=IM<b6HWSc7OT#Y(K-]TPJNbeFY)XUF8Ef:e0+Ee.JJPUQHJeG
U+#(XHe;+Q.a(_JUAP4_:ST;GR=HZYDT>IHST?K&L7P7GCZ:W2fa489UaB8a,;8H
L()N<-+67+Q:/OJ_.4NCR6TfZMXU<W4Z=U^b&6Q.&D+[.,O\;\G@fILI)d4HW93^
CIQ0BcKfAI^)^9COGaJN]XMZ-A4c64gW\&(]K;R&4/8/bT:CX]A,<;>->2M_H<Q#
QLbP]afb7#>HM^DT\8X?P,;C#D^Q5>VE165O]RI]#D_41J.&QO4M+YJ(+YN<\>D)
>Sf&G39ag^OAW:f?3f380CU[P0)9b=ZH2PN(_R0-6d-@RHB=J&=:\8UZNDY>EgSf
#g;5D1]H6A[8E^.B),RAG^b#DYeE5;FF(-65E_42,]6OFcA\HT691C2W<d@ET6Lb
CIaMLNAfZMV9Vf9GRR[00=]b\=Z@J6&aD,78cLF]]U=b6@f.G3;JDY2P47;]Y4K,
9,B5WU[NP(M7=CEV^=+T.B&++CO6(LEe?YB.9&3&Y@;GeB+J9(gIS&d/[7IM2]I4
ILgUL&O]\Aed:WF#4_=.c^208H)EUPA?=J0VU.8#CRZ/K,J13,FDd51AfV^?D79W
4QDH>(-UHZLIP1OK4J,>V^33/[5&RJ+eLS4)a0g^M\3PJRAOGXH2HeeM:#=Z?Pc.
9>8[?=+2\#;4YeL7-U#(b).;Jg28PTf1N;gH[(eS\STe:HKK+fK2RY64]d&5:d)b
/(e\^e#:fcT:@O\:XO+5;M)Xe^ET=)&+gZ<:O7;CH/Q^LBf#T;,7LQ]JP&c2f1GU
<gY_-J.HcSK3&C7OcWbC:e^:\WM2e\H9I2LYN2=RDJASeBCZ3&@]AgM:^3ZK7FAa
2gY27([51Y.@)g7&d&O7(Yc^;BW_1=A7cC_=ANF-RBFP)2U)4bKS3B0,>VG3S=6J
&B6AW;5:-eQ3@,?dKYYLM\7A\eI?@dEd3P:GGH+#E)PD_a4R^/b&&0@Q=TSW\_\^
T.+6-\cc71,-N?459HQ7<DIW&N8?+>e]eZXf4UcX+X5g4JJ\\OePH(5#8C:79Y:0
E[cLBL1b-V/1Q[>6;D5H:2A/;8\NQ&BS_^Sf^7dS=^DF-KA4X>Q2J.--IPZ5(Z6]
&V2Fg1B]bBVZ:RH6ITQ_]GLIVa=@]e<^;cPb6GJL-])6f1gOf2DdJ_)/bL6^7^_O
F#78^9V-U[5RU46EP3]NbdEb/KH\<YK[/HZ:(:Y?)NfA4A1faP1E/b4>7dAA:M-P
\e54FRON/-<dcZ8_TGV5R?^GA9;KJ#RY?g\OP?,c0T0c26DYcUIC48&Y/CA:;0@V
=1P\)gJ@)I(Gd]E9//REL+80@2O)-K.43\?7Jb)/NeGWN;ON#B1X79.>]+)P:)+0
#,O451fH=gLN@G8?3M4:)N&77V9:9@=B-V(K^PX@FU:1_:cSdSf33g/^VY_W7:fM
eH^4+;9)@<PXbAPfeEG9c7&C>#SL&RgQfMd)_CNY\b]_R-K#X;_=:G=Xc:^;]GHI
Y8[/O=S^3Ea_^N>79YQ[J+:D#@c_6IO4MB#1bHACSD;EG,_69#a-\Ze#V[RX8fg?
^\c18/Ud.=3;/1;UT[W7Y<+6P7/VH[S3(HL_31>SN;3JM]>\LIGb\=e<6HBO8DJD
+XgKXbRfT.Y&CbVFXLUd4)Qb@Q;:1E[EU42+O;OO+MXe_HZTY7.\F?,^0f^XdAKC
KOOY;+CTNeRC1L+4:LQ4_]T(9bT]:<Q8([U5V1GP>N2]#4WSWUc,AW6X^5N1K6#1
dcG-8?P?d9@=[,eP)G8a?O3KFA8/__f\5f<a5[e^5bF[b\=7+K5U+D3)UVgGBZ#;
]O(,W(H1<#^Ne#6IKI+MI9/g?aTGKUeX5/GCV/@;gcg,U./3(GUR:D)Zc(eT-\6H
)]1)&BI.f>;HM5M,J\1L++&[C5JUcdY&A2L)5<H4?c4YeZ5&[RRB0SS;,&.BVcM+
T^cRb\<^eO#;b4[WK[WVT-^.d,HPYb::^,ca57(-2^I.;:.T\.^WaO;0DH<<dK_>
(\IDW^<=F^_6,^QGgF,[39I@E6)dN5=:(5OLH2^G<SbL]U4A1RG1F]3<S-Ag64NQ
D8@SXc9Tbc70U5G:O^O>Y;g@;YDE-X[>WS4EB,UVS<.0+J)H-#G+gceI9K6XUb[:
\+)#&WEL)7[^9W?dV(5#JALaQ==Q65#>:IIQ>DZXMNX;\F]57;51WBM7NS[?fc.:
VCQa]\WH<)1QD^NAY+ARI=A;L:EMeP,<_5ZCc607:GTdLK(G],_8^^-PB><FDLE<
EDa5)H8H,H#^^^R3LZ^af5GE7d=Ne&W[NPS4]e4AdgG\?<BD4RfP1_9W8@@VCA3J
7CJ>aL.>dULXf#)0W55/e&GREEOY^KS@&2&NA_38bDXLL><W4/+UMAV(VF.ad)5N
F;Wc,:]_.D53430MZ)^AY?Q[,&WgZ3XdGB+gXVN4@Q=dbM9K9I-T1,Z;Y8MF_;WZ
V0_L+&WG=E0JPVJM?GID56e8-EO#ae91RKE=HPS&c)B@9N&>5.X4AO)0Fe1EA8/F
<]X;NVP5S3[E\0F5d)4G&6MG3+4L^[K0I:Wf);1DWIS7,>;fN^&AUGe?bA>#EV_)
RA4cW5f>Q,gG5MIUd(@H4Zbdf+7XVbdP3Z&e[WHf9AIAGdB)+WD[<KNdM6+20KaR
6/U5BF#>R/Z_bag<3Je(#T>2RCVL-a[4D(XP^=+MSH0(JcE]e@+.Q8#VYB_.8g):
WCWC9<TOW)1O7E4>1G4K)4PJ31<TC.&AJc7]U<F4RW^D?/FUJ_SZ\)0#>E,cb<1[
7Q5P-NBbLJO;@]>CM4Y:9N(?06>91G:D5D]]fd3/=&Ed+.bQ)0A57>/)DD63V/[b
E8-1Y&BcOe:.d1,L=<1XaPV8?GNL>]Dd,,Y:0[6\JHZIaLQ^/_RGT9g8d_+?NPN3
L/VgO[J1eFJ9S8F5JXS;?E?5<JH<1XL.ZZD2WE\VSAKLCZJJc6>KaTFJ7XG7.[\6
8KAS173^BP@QgWC;VPT?><G<W/#EgINA4BNLZI1H19Y<HM9D@&eXSN91N&LJP:g+
ZZJK<7@RA;c<FYeK#1UL[Z?&+GZ1g)Y[RWSWgaeF]ZVF0=KL3RP-B+M;&d,Tc?e9
\6NPeHF,N57d[4FKNC^WA^YMM8R7B7(]8>(f=O#D]e-I?V.b7643P7MK3O1>V.+I
37cM20TJ85-P9.LY(BKB1[RI.[3W\EM2[Y4XUV/b):O,aM1&7UPKU;54UVL?4J9g
8f2PFNS@U<IMWAeN;E^Yd,7(e]LAR\>eRcHE5#9:(&YU6<>4;)@9T0&>J5DJJ\02
_Of#NC<W+C;c_AMFQX.64#+Of^:4JC+0^VNBVc:^A8IBP8d)A<+fbf5XSO/_GUIA
&WV:.C9@NW9b\JK+.0F=9aB-/,JgG9N6FDEgO#VU#LX_3]DMTgLg0CJ+JUW-b\Ag
-_[]&XA>eC9Kd8=,ZSL6PMU:D?:K59U+I^X=HXD)>CRbK+L8B901MO<>,5X0IFV=
N>DXU_+B<8Z55SXZ1+@;@deJ.\[1U5A<MEB,Ac^[94>?)K0deXSU6ff,g+,RF_d]
ESU6YfUO#CZC@N:SM<8P?VB0+LY__1_Ab3G)Q)U)6a\1X^^.FJKC9e2(XIg6&0Ig
P#P_A1T0B<_C8M;dR1XRY,OM+BW7U4NN;K0?8O??-5H)@8K7RbCSAfC+H4G\R&)W
#e)T;JI60)8d>+4G76T[LO9ZE+0b.+_.bMN^Q+YV\Tg&6MOLU:EG-Q@SDR3+J(AB
d<9f^gb;aB.W2G,?dB.:JE,YF)c0+WeJ.2(D1N=#0?:EO\(LA0K4RM&Cb?)bW69R
0?BKR<9K./7ITL?>PE;9J@J<eT8.Fa-T4P2.\W.V+UQZY?AH1Y2_]M+NYBW_>;L/
+c>.&ORd\Q[f:8g\74?HN=#-d8Ea?]IW3\EfQa;L7gD9C0,^OB5g9Agd)INLIg:?
d7//I/:Zb)(de3RKdXTOWQ1ID]SG4&O^DYIY<-AcdAC=f<fR#F=/TEKS=BNH^@..
0?]I49cL1C[+7_49I-+H[6,GH>NG)=QeO,Md[DNBPM2?.DT#V-2)WT#=,=>LK8(4
I6&UWa\UU4Le#6(K^cdV)aUY]dK>\[M_?=\R7-_30B[..^C,@]K^E[ICDGI:#HJ;
787Z;f8Y_d-R&72/_L_K7g@\5SQ48CTgY\J,6Ye0^T94#25dU4&G3.M:<KV,[@UU
,\3[ZCHHWAb6_/S_Z/ZBYFFQUH(TX2LGWD+9@W-[=@96_K)62)SH;0KXRe[d]c:G
F/&R6a+^;JO>Z@K1JQf6>Y5=JGNA(4)#Cg2G2=D#b1R]V&5G?));_GV<PA:]JEeP
VNU<6.JP&^<5CD;O^P6IP1?O9ZBFSEGN>>eJUeM76NE-O&3bgW1Q3G4P/4_.1J=1
.C-=(D\GMD6D2OXB4[;#R0Q@bd5<PXGI:&1KDEK^IJ1YgO=1K7R7)eNMMRcT>E#7
2YOO3<F6I#Rf_+&@X\=ffU(;A;<f54IT4VT1NB(BA.b9VEK(_7Fb3VdN#9YU4>R#
cWXAd#5ZHeKD_HC((5]AIfZZ.M]Q(QQND,>+5.e735JB7Bd0XY>gbH4YF\<,5(Bc
XV98N5[O6-(.H+:@>\M[_L1Nd?M<5U6E\4aYIW_?^/]_#XJT?XV2#B(4G+EL]c5d
)c#2/D(gCTZ8FMFL58+e=3]&#Q,14L:6U2M\8^W=S)Z^A0.,N5bM]FDX>-_1W8YM
fD0J+FQ3gGS>]TPS-K5RCbI[&53>BeGHKO\5D#48[af-][9GC+7@S,\IMKNd(30S
?-KA6WK1#Ib/,Gbg(KF<G/Q32&BYKf(+GW1[7E<?;M)1IO1\M:eF4?-bE41&f=7G
2f7BULH5)&60@=Cc.SQ1;5O&#Z_d;,:T0-&M<+^KQ<NILH08O(Ag#HRKfdLAcTL#
2P>+HW5EERK?GJ9MY1;1E1TRD._f/fRBO>7fcgVNTU44HKKV(ZFeaCM7T2=fDWQM
HA?7g:CK]f],S?QV5@ZSI+?MJ5cY#H#ST0Db=]0^+;4=_]/ZN25<^>>+&dZ[YOg#
=^=(-&&M:K6d<DJX9;@?c\_F?^)I0P/.AgK<.MKHKP6>X;4;.][fW8R;>eXM:>aI
[Z-]Q0FVC9O_>+\A]W5IF2_Ha5gBQFW.a5P#G5?JHJJ4FeKQJISS/IA<>Pe2ZS#?
\9KXH8+IbG9PXKQVAcWIR^8#)g7W3IGg?=W.67&A6NL&WNPgTbgDVY5+J:g52feK
,;=I5W0Vd7PN8L@(Z\RQNC9#\1#C1,We6@@QI[gJ;:96OGg,AC/_X4N=J65[\ae0
0cU[N/&\Ag+X7fgR\P@\+0CHg38T[,X;,EUFPB.7<7,Q(GK3)#WZ&1/DO1TLG](f
-#Gb3,9@O>X,(JZ+B2MadTN\;f/D\\O?;P&E86<Xd887fd,Y9+>+&;O0_R50RGCA
&/V\57e;N&^XECXg_:6[+&:UH9^9C;H&LX@]JIPG>O1FbNN@LIN_R6F#4J=VSTa\
8eAP^Y\I#)Q/LIGHOKK=QQ6E.50LZ,4ZS&ZD6TCeZ\b4](JB)^@GB.?AT4VdEG=f
TOHJP[80/=/B<\@ab5-[?A]IH;NDN:Q3<QCQG2H-fI]aKLGC5&;\WG.DAFVS,42_
<b124U;G4;->2/Vb+A&U:#C/a]f@]0J9QE@#J1T;#]K57D2XU0T>,0=cC8FLLFC2
H>2MF0e3WaM2Z-ML9ARON2@K5=RK.]ff(28I>Lb=];D5.5C@QXS=gXVGKZAQ_^G=
Z#3Y,RNYE8A-Z3RA@&=Y@.H3<>A)CDV?Y2J(Le0LC?;J]f7CRgQ-g;)6-\^3]Q,T
A)(6MdOD6B4K8^+>8RYQKE1S-:J?^M8B,@ZRbRLF+f@]BY(0-cS>SJf1\/9W#X,T
S(&^]>aXXgA7T)9a,EZ@5Z#F-LVYB/)2E2()RJ/KDYMD_G>RP#fYQXPSfLDb&BXQ
8GCb5N4WQ^bPA62YU)D^I^ET-\?^A1T&^E)O>=8;U#/@D7O,T2Y0<PCPM2<<E_C[
AD,:)&8A/W#@-bc/K2g>^aQ8)JabH.E;.HB9AP[Qd2d\8ZfSK&[X_>MY0D#&1Sb_
^1(gEcHJ]MA/4;WVeB>4Ya<-WG,=AeY9X<U^/@b.+Def@BU/UTD0:ST(b60>d2FU
OU>Agd[P.>VDMe7^\SPA25+TS312bD>+H8E5/_)OVLdW(0BQ>F^)58DW9SD[&,0&
C-+6W/.S2g[b8dR>JNKT<JEMP9g/3\/bPa;78>F\2e?SG^._VW0g,2<b5)=ZHY,]
/Og8FS9D<DN)BJ-:1[(ZGGe?:_PW.9gLOJZdBF+3f_<6d_NS6JEbN)8=fGKNGI7O
F[?_Y@P-&U.WA[5PdV+1a6&fUgX);8/8db<:cATE\&_K3&^IM33)35Q<.R5L):D^
=A(BXQSNVe<8Z3^0OMIVQ/J4)N00e_\)M[J[K#;1MRXUE2^Q5f]0OR,<G4>Y)2gg
2.YN9VUQGF^7[FIW9E.G^Le,MPXT,_dBCCFY5:4eB1V4,)QeOcXHJ[\,/\T[R(14
#eQ5a6e_B[QO36)?PF&SXXXM0F,,AP35QE=O1JV/WL/5GEg)YYBd<DJ_MFe5Q4.B
/<DCSDC2,W;KfIO)PG2a&5@JfC45B#DKf137M:K,d]T)fdY5RcOVDYdXE+XIHX7R
X4AD\-I-.93-;I_3gBY?,YWT&Rg0Ka[JcI2GG.M@c5M9(JN/d68MJf?1]2G=6R1V
c@0ffS8fGY,CZc4+M?]Ye4[CE1]WOXTQf4?^>;[^8=XKC-2SS\(RI9&fgDR<RXDD
Fa4UA\5dU9+De&d;7d<18Sc.LU=eH5Q#HN3bODUC>GJ,SL(2+[^+e.)(\_D9T;X5
NJRcMQD#;_G.72)888-b>[cE\.#Z:=-^[-BI0g+KF-G87AI6@7KeaR03c[b6X-d+
:AId6f3:D]SK3e8]@468VPd&/:30\AW2Y@d,<1Tf[3cQ<MM6T+63Fb.KGg+UA(2>
-)8IY9\:HQAB>C=5=QTdGb-5XGR=GP&+EO_.7&?b.1Z5@U#(#>2<a&_T(GG]Z33J
T]KN>GEY5<4,]7dULVTZ)HJfC,5gB-5O85I2Q.HG+gEI,)B\8Y43W^QGg3@<C/bG
KFJ)c)A\2.#D47EU-AWFC/J)6<_CJ:OG,.g?L<O]-a->CV6FJe_U-3),-\eBBB3T
?(S]@N1afTEa\+A9]1U=#K]Q<?4WZTPdHH_^VBX;Z(A.A2?2@7Og_PcFLO&_cBXI
f[6WS9NQJ@+Q)X.L#[cfXEYQIE_^DYZcPUc1HS@/BSYK5fS>I.1J:X#FYg_HZ6bd
4_VVaB.(NdEER\)Z=^./eBA]CcG)_f+OT.@G#a_J+>-+8[HD2#0e8?LZAF.-I2cM
B7Nb&TOa(&Q:L,f:)I;Ebg9f6>e=]/EHAQda\Z]?OCNJQOGfbV<XX<d0DZLfJf0)
3Z4W#F#T5a1dH.=57/^B(PM_g7I/QgceQTCMdC/EK_74WA(bGJKR+5-<XHJMReID
\THHNB8QHPZ_.Y72W-I=Xb(?M&NaD#ZQC/@VJ^W,bV.c3Sb6Qfc#d4PL[;2ZP)H.
UD&Q-&b7a&QH],[^:@DTO;ZW7)\2=D^@RW62(Hg-3JRdB(^TP-YWSW);_MIC;2>=
Wba-Z]2#aS1[(Ec,Rb:F/=JJ2(W^_^R8.KVAM<Jbf\\BOZL9\9;/aPAa6<CT[C=U
La>02(bZ.e>[9P2bZWc6bJ4XdPI3^\5@BQ#5[=[A+JW0A_C&B@MAZ@EJT/^IHbQb
G7((b^;PIH(V[Mac?OE&VQ4?IXg&&,,GLY0P48N2W#a9>:G_+-C/gIOC8LfN(H9c
b1Y=2L0FQ=R0N_J,E??K[#62FX5>e?]>G9T.3&?X29)H&;8N?U/eT_3L>-QE7W)Q
X##UU6MV-J/@ZC:E1EUK:D<9V<;c@5OHOgY:>W,0>O#8#TS,&FWK_/c?>bFPM:B_
]ERfHFG6dCZ1:e:/=T_ZZPFT^D[+0O4+/<+];2\N8CF6d(E5])U;^0;ZX1SE&)35
R>7BL)2d7G\>U1=8&4/N)3Je6?b[GU(B82VedbS0fRG\AJdGA(?RH:?+>YE7,FS@
?PSN=1>EQe9eNcKB><cF::2=ALQ(IE^=?\CVRV>H29bH7eAcBN.TJ)U3710SaZZW
M3#N8W<VEdQc75Z1efGP(C13N5Q@71NHb]O?6IJ^.?.2<WW_N3aBN>Xd?D1RPTP1
@0XDG2>A:F@YIg^>]P]81-e\=+g:#T9J?f19]^^?+]=[+,ADND@4G1N3aI]0(W?.
f2_9A4\P64XEWd8[Y#CKa3]62Y^@9aUIFaCP40S86I)C_ZX]E<WL<(d,+L.\Hb@M
D^?;H0fBGJB45W]M]?+9;,F8.g5.Z^NRBYOVTbC4Q(>BF9>5b,AE8,DdM];0T#V2
6+EW_[JJY))_M;e3B[@T,E2=6QYPHQTP^EdD+X;C,G18/2@3a>f+UZf0YX/f.>g&
CBf0<[H^B3d&_===CYRASJ4b3C2MaP;SU8eW,<RP[-U@#4I+])GKO<75<GT8TEcf
,#+M5J+\^TM6/X;E2X,W_V;QAO[OD?)OUDEbK,=KPf_4Y+NaQIUgb-:]HL5-U&4G
Xc8a-NFZN\B[]L>7^Xe.ZPdc#/>e\a.6KbP<&3/]])8gY,-1ZgUg1WLJ>PDEA^X7
@O,?LN\04cZK59<\)ag91[B.8[(C5.:)MP0cKJAXSK-JL(AF;a@3]Ib07M?G(c7M
,8ae\(36eSGIS<7f)?&0f9GH-.f\d3N3W;RX,Y@aB(Lf0ETSD:NTgK3Lb7H++>_N
Wf2_6UWV+\>9M])3Eg?_XN#/R8=158+32[<^NX=C[:3F[[,(ee.S_c2#g22=LM.>
DfRbgM[=LXb/YHH<gT#6C(Z:@f_00SGK\D;Gfg9?FIc<_e.4&]#)e[#d;YI?f?R<
EZ)+-[eZf]T=@BPWPX3]Xb7a(SH(\PN35?E&9V^?W4ZJ_XOPV[CY_WD@^.11ZG/6
E_?=a5^4U?_e\DU3[_M]&bXRY2M+dZ-LW2S+F:P&S(R(>8A7E7AHES=+3_5>=#d#
M0Y=O)U]e]M>N,1f6a;?1g=B#1GKLC_>[@\gGE:@D?T4^f,N^H/B6U6V++E;U_L5
L;:]fV<A-RN6^6P)cO-Q#J6gGb04V\FC49A3<^3AD5.#BM4JNO-:#LK(f[Nf1L8<
2aAM,Xd^9K=2a5;R.&Zg]FB=N;UGeD)@&AD3\.Ye)3JGU=f]]+c,,X]FdN?AOMGQ
7YO<NIEb?@EcF\-,?PL&[K1=@QG@d_Re5D10EB#V[H7FdWR(GJ72?[T.QM0#GDf5
#4WMYQLg=gPLdZZM=ecSB@_EX--Z93CZW#BP0dT]<XW[Q#Wa8?A;?eaC(L#[UE,c
#X?f6>bbBV)DU87B,1RCX1841Z7V0C3YL]N[M/\PU+VTQ^_50^<J33(afBIH1NY^
RH=DaSRe\e+c>>9[Q(f4=a;&),cE.dGO(T772^e&?9=RL)-K+)XCPNRe>.2aL0=I
=.6Y\Rb42QCI>Q]9BBWE&QeT1Zf.WR57OWT),R7O5N2/WdZJW9P,0KG?G2,G4KC<
4&6&R\)gT+??XWKXDaC=0CbB+^a.#O_^GWFT->F;Oa[(G0Ze+QfR-eBeUg[_J?fP
20\U/N9\ZV_::/.:I<EED5/E;_L8(SfM)L;8IC32V&0\V1U/MFBgD:gSadMJOQ13
&<+GOI]K/2)^[[\[[OU:))cL)USR;<4:N\INML0\CE7M1<&U.8IN@gV<Db\SY+>0
3###R7@M;E@dJ-LRd4a/Q?W184/]D8_(._?WG17LUM.I0LXPFIEdPW3A2B]#O41P
Rd90I>9\bOV#a.@_1U,Q=RUPZGU[<IM4F+1<<3WY]P=ReCTY0GTgERW:aO)@V^/<
@ggFDNK?O5ddP#6B;#Hf9dSe88JTc3.EWNIQ;KUDVe=4.F(Y6dcT#,[eZa/?15UL
f2PcT8<-H3c83=PPO>V+:]=#1/.XGN-O)?KL\KYfTRKbT:ba9+JQbN]JH^ZTEf?F
O_4K4Wf>-)g3Q4^d08\,;d6].G+.[;a<;OH#_UC2Ra0ABR,H;<)62B.S8TQJQcJ/
<g?M^O-.]=-.T/B@b775D0SJ-PW/WJAH27Yf7IFE[;XHf/A6=Ca)>6XV5C@,g9e^
;?2DC^]6(Q>e6><c(GF;N<(RDK@b+RMH76CT/=]]U,9XOT1-QGG=PREJ.J;/Q)9F
140Af1+[(AUP66#DdeUDO:[@H/6:(?2@X;M7(N7LgdD\7eU/0F?e1NFL,\GZJ/Q>
g8&4;KZGGJ_aa(P4ID)]5Cf(f>DII?6-\7#(#DB3[<fHC<L4I<T?ZUgQR4P_M^WP
ABJK:50?@H+6Y7Xg08gTa^R40\W>SW-14]Z?DXO2d3,&deZOdE2\.ZQ1g@b=b)8Z
]J4=9FUQZYd3N+4\Z1,Q3QEVAU9WJK_3\PR.K4[Of\#?<KgZQ13;ZH[2EXAXOQbY
I(I1HdMC8;U8bMP7R=Tcg..dDSVK&P@>=/aT3>aPE@=R5&;CM+S]=EI5[FEMC#VE
FU<[MQW>5JUfVFY:&&5P9)a+8N#]1H)9&K)[O&EX)&>5W.H+dXe93g_,NJfa(I[<
.QN_e<9cb9?+R](\#LJXY/3(-He@Q;0C#1@2&B<IUOJ8B^4>_HU?TP\[53N6=_WY
BQeFC8?MF:,FEPA1\1)QbQ?X-,8]93<T4N5J0H\,+._(P36N4W3_A/Xg1/QbQR(g
cXDQN\J<fN?0#5QIP[bLE5W.O)B2D:NW1=Q[Y99AC4;#[d5^?Weg#7eJCKJ@A?Y,
C7cW-VDE[1TMbb3;U7.FD03M#T,]QgQUUEB-N;3UO\BaP@]S+1J1+J2-CL/c5>6T
?cU\@&B]5H#:eH4&Q3)8@UYgM6Wd_ZIU0.ZW]a^6W.f6II3f+ba:WQN#a5K/eJ7S
2N3fP?\#[6BY#a(DFeF.LJ_])S_=QFL(;E>@Y^561X7Eb.4Cb4.S14e4_-CVK,1N
&;1&^K2SOW&G<I=Y:LBc0(I9=K7/]9-:>X\V7@MF==]7W_&C\0THQ)^N_M3TaOR4
F?T0[7a_B<cc1P=cM85gb1QRGf.JFF\Q[6(<J<1S?S-\H];1X+DJH]S#\cD@I/(J
f<=BABYTV+#1d#c48]g<c9FP^g_J<fQ27NGX9_+/&GXg-MAR/,X+#FDP5RHWc.b9
A3CUR?)3/PSgOc)4Z\OLB]IZaX9JBO>Z_OJ)JS.0/^ZRe^F[PaC?P<ZBFc/4MNFH
QYcHW94&)f3GIGW+N?9Q(-C96S9Ae7D>B3->Id1DfQL,\A]/1GCVFQ2>WZBVRCLI
3E^]N?Q4&52A_)_/NB4ZY#^@2;fYY37_Aa^IbRWAee?Q,<f1@?=]J\gZNDRA)9.<
8U2\UY(,YPTP_UPNb?+?O)F1f_\RAB+K.(aYPM#=a\N)G&QOJT1[<W([>\Q<9H_@
/B&>O-D\..53O=4NWAG]6P5SI.Yd1G3FccKbSS#24cC,XJQ=d0.[WV9F2f0aSUFA
^S<T1\<)GI4)@9e3YZJD=YI4ANCZFZ>+7RSTI\Q>Ta)7Z<P7Eb=;[W\?//J+;?&2
bANBP(<X[B?#HYR7.,V+f,@CN.=7_REVL-dB2#1d4;EE3#fPGK5ZVDBb:>[e\G=F
)UR>,.:NXc4KEP#L:;1DL++/aVL7&YVOD:97A9QO_T7N]2BX79XNa.Q(J/ZN7107
6\WK@4N]969+fIUgY_Y]d.L5#PgN24S)\9NMSe88D]Z/6A;?RTS)@bdQNZBNb@K>
QD8Yd81bC8;afRA60@+FD7YPfV1.CcW\:--\@)FS9:2J>CZ\g>aY[b\ASJ^Sc(O\
Q&YP=e;?1>+1/=C+[[?_((P=]cf.\X=S=+JV\?3cNgCQAM#g?:Z,g&XQOYB-JI_D
)W[0T)Fd_=a#GfA;f-b23>N(a&./e0gG_[3>aK<^/ZX#IaGBT]/@OQ34@<2J))A2
#S0#Z]fZ_c<BXLTX8\OYFF._+>NN7332MLHXaHWCHNO@OW9a,bM;EF.fZ9V<T>;.
=48<7LEGYOHL>)&8[CBAZ<:6+^+ZI@AE:#_T=_37>6Q3)>.@,T:f6>O=P-3NYIDT
3NAODAaGR1_YDL)/K.PB\N04S,L^Ta,S&Q]aA)e1:Gg&N:1@2L.&QR/&CT846W6b
LI&MK8[XO^9P@LAG?RO[J.QG))0]1c0F<+c@]:THHQ7TJ/XM,3;>N:B&24/JBg/@
C0McFMO]ZV^>Ad+_-CV^&FXT>cbB0bB[/1333_->(:,]P=C=QA2VHB8[=]-3XK;W
7=1&eWCfNY,79e=4(dZ^I,N#JZ^L.2fHD-48-^D#Oc,TNAQ_X4+T((1E\\C=J5OJ
./.Qg.6MSXPK;E^+?dK#7^JY,RWYAZ?R>(+UA>g:a72WZ(70aJ3\<b09geMSCST@
OV_OaNP4b7>5T9RJSG8^=QU-9AWIHB(4&]6YO/L8HEa5\M<\2aY4YTYMMZ2H:(3f
W_=SA=EGI)1,FS)dLKB)]A@8GB2T:e[ES9LN]F3)@MCGGaMRR^GHJP^]ddcH5:)=
)O/:GQ8R1/6MNPK_7g#>SN4.Ue:dUVC@]I5?H#8U5&&e1+>XH99Jf>&,,LLXB2[,
HKC1UVVf+6I\D(R7CL6@^K492K3>;WP.Q4Q;A,<^S5S7=DLK\0)HXCNS>bR1#g.2
KNC-\aZd7EJM_a7=@b:KeeI-<]C(R?9\/368aCddDNVd?Q]&#a<0>8Ag.3bHE6^N
FH:M04VM6:;^XD^?C=RH,H_d;U7;A1EL94M]6>//AF4I/+5+Ub+T[R:7#UU;M1CJ
-?g_3)OPK]#Pf<-.cZAXJ?EBNed3SfV2V04c/?OQE9=YP.C<,ReC50YO:=IbDLX5
e<YT9GQJ_E>Tf>+IZZX3+LC_aP:YMP:8SUcPDFO7F6F[&<L&W26+@_<;/4.W9L7K
-dQSf]0@Nf(Fc[^81J2;W@#_^8;85QVS:B5+PTM0.JJ(?Uc;K7^J)Of49=T-MCCg
V.V5[.#;OHW\?4dA;?BG[)2PHaL@30N6#IA9A]FHE##Y9KG)CJ0#:V6@aZRPH[[_
>S4H,d/VFcD.,,S1[&SD]I&T657aU]3)Z7XQceBdDR[N9gcS&VSH^E7N53(4L<PO
VAD4T8F@N?ac[4[M@JW8K]T:4+<BETMRIJHR,<Q=UIXgb<dI=0^6Td?c4QDM60L7
03g0Y.M0I0gS3+=(4VDbEGEQIbJNGa-=\O6<a)/1^#H4S[:6:E0.S0L1fFBR^#5_
HPZ@g.KPSX<_A690.[Hf4e=9f7006?(6+0:cADP=J85,0d@L>:QJ/Pd#DK\0M9b_
c1a1#_>VZLg,N2ZgVAC(dHPDI]G;ef#LX5UPOJG6aYEC3f5U=N<;@a.HOQ_,.8>M
W@Q4b&0c,F#-7=EP2VF5f6\VH3)P52BDAd]3GE07MN:]/0:W-e/0C\VVc5J4ebB\
LS]1af2.A4+I,<Q,Z>Od(g[;63^4:PDEYI(OXLX0HJP8>]Eb(O678Ga^[5fEQG#Y
QEFe(:[M8b_#TM]DGT:=bT(Z?AZa+DJ419Rf5N>;EOO(=_&O=2EMU.10BeG]-XKP
E708Y[^1;/40W+VV\Q^]?3>52a<OZNf^3)4B6Ff:\M:6f3BW#)-M4YJA<05)AI+g
QT?(7Y9?_3IWPOO,.E4QB2KEJdVTfE23-(8F,-D5D/g;2SFc^MRD3S;aSgKN)ec)
9,d@ggLQe8.c,05gYLTa>>4I81J3QQS^=_1U/7ffUPKT&=GV^--7T.dMY554A5U)
_N;SN96SF++Acd,TWMJPg^HW6@,5W\F1PbB^&HCP&>F<G&[/0^GH7PV&/33FN7?8
0KG,.d5I6.H.CH[E2[[K\:.AQIV0aO?YPR?&+\_[I01c-TWMZMAUDF-c]O..&A-g
7\,P^eC?J7IZ&9WCS@O6Bd([@;:g&4-5--gdaJJ2aOD=ag6R\B&P^3M3#RD))_b\
,RR54X4fE8[]N3QM-34e)Z+U_HI+9_Y9>a\FQG08&@RK-N<KLZ0MB\U2=;cZ8Vcf
ZZMCGc#5e1CH30gUL;F(7d^UVH7e;,.Wb_#LdY)XHN?7RN-16GE:2OY>J:@,Ifa(
>;I#a/X&G/HC)]Z(J89Zd@_,(Gc(+0U+aU-E3U#>1_e87KZP./1HE;JVd5PQ_ACA
,JK,N,IY=J+S?IQdZg#L9V1VZ:(^C68ROTKW]5FgUL7HC]_RH9VBZ8gDf0>#(GD_
H_U?W_,XU@/J\:<A-.]<@OO52\\Pc_&^b>gS;=O0,_6c_eL2)U;fW7@PWd1bDJEM
,?),Q3)117>4;AG=CIAME;)6ETWL\]NO>gc3VaJ0KA3X]^)YLG4(c@7f:QQ6K6[\
<:6ZWQ_R?ZQK8;01\OBZa@ZY??UQ30+052d##;e),/e:Jb?3OVEDRb+AcH+HWd/(
4/4aLNDTVRH^5f13bA1<2GSB\HAc8H7bL45)>Eb2-4U#4G2L[&Z,/39T^MNb+=?b
R=D(e\6)@T\MfO]:CM;KCV(V4VK:]:]F^6dK;A.VCS=S0RRH:dGPbdeA\5IdH2X\
BbB0@Ga^D,?J4,)7N#4cXXD]Z<N,XWNAMZN26V_:ZZE5/^D]^4@@R61/0\SO5F+#
@[?GRIZ+87&=K^MS7X=/<<4gQK5LZd@gc(H2RNL+,)WFNb14Z8S0S)<_Z[Rf]&Z;
A[6@N&>CX=AB>4(V2(0dbIbWY(]N1SEYc_/+Z@<daNHHQQf_^V5YZ6PTPE?\0_Vc
f-7Q=5/\3O]@N+G6P9B#1P^6T1TB3T=dAQ9,42=HCAWdIQcF\P,XEe<?P-6WE]ZL
-HMS)cdQ4.G)Kg]bB0M6TCbW;-JVXP&Of6V(SC5(?gD<L.:eB,ODTd4Y<2H2SB6,
T/G8[LR?S)BcUU5B[RKK9a?1K;@A(g&RBKUV\4KY_W-?^EU(-e9-+?.fA6F\gaM;
dA+8aZ=,>.:O-bMT(87RI\JKK.238H,9a.P6EWLWab(S.HML-a5D>S6D:+7&/TE[
EVV]YcMTEOTG&3De/gM6R:?#I/MNPE+X1gf__IVVLUY58Ya.,EI1].#aLX.4M[g_
0:]2>.be/RW3UR+:XRO&1AQE8.^g9g[2K\<1gYL6=-OdZa5\(6#:_,F/9Z5F?WN6
2]@cBeJ0B/8G?gWUeb5VccKcS2\2A6H5XR6:5EMLJPSW.UZ;<-UJC;ZKHOQS5/7?
(:XG2C[\Qc;W+f@>:gMH_#2_@Z0IS#TRYEeHDP>WY2_3QF&aIa<]F56E1<CZ:9D3
/<b6\3E4eSZ.Z69J_SF2OdHA@)&WHeGcg)Qc,748XUT#Z>e?-8_5eYJ<S^8d4.\8
;4K>L83U23=GQX2\a.J3;KL743Y#WOR7-N;=fS7PL@[;/bgS5(_g]<-2KQ&NdT,L
\3Y\/.I&YRL0Z^)_TI?:.Abf4fRY\_0F7:Qc46D)1SP/\&\A3]W8V[2_TJ^C.:2H
dJ46HE[=RYVYHO2=/4OUQI=WNOI/\TOY+V.)B1#O=N=g/Q.HfeHE?(.8>#FQdI,7
b10:AbM;_2:,R?2ZGHH=#G2]9HIWdW5R#>QUeB(?WH=(J&+T[_DgCR-fSC(]Y+/0
Nf[JHT)\cE=VO_:O,aS6J2FFO3ZR_I8H,0b^b&6Ug&[c4+c<C>K:aNdP0\S/La3<
P\8@[.M+O#575V.]f58gS),ef&2IVL+:23V;5LgKVfbK=K>1[/e=ST5R;7?<U,:_
AJSI^^H<]A.-&]VDT76GTQ^\?Y02UDgVJWC]>M\>I(?CR<(\CgY,)B9I(X<>BS^e
]PC3MYcHH??gW)/8YU[VR/(Wa@93aWUYTWd[Z10Ndg&I3/&FA>QH]DI&\9+QY\]-
CaIQBWg2DKP4)bd6#09TbLV0C<0XGDb7\ZRM85T8>?c\B6YVPfQH5FP8H/8L@ee1
YP1f=<_6:L:#VYR0EZPL4bS1UX]@WX822+]V&Vb83_gRZ/O)SV7<U4X;W+6O]1^>
G>0ega8V:RN/1R(d95K+AIVf<U<XgEI[KPaeESf4I@KMg<80:#D:dRL:-FgMY)L.
J=.41C5S(E[:Bb^>&:c(-V6g;,J24LAHU[R+#4aHE^Q+g9NeF,PaAQL04=Y.+O41
\7=7;Vf:MdXfbd=]+D+/96SP>P]NbC><JN\&A#2_T^LcZU3LLaB()VE4@b[aV1Ab
:>M_VW/CZ_8CD+9EV7[0_&Y>WeG9Qe@5178_dP0YFBJAE>cYC(5bOMRBL-4ZNQ6_
51H4LGR9_]U48c<]OJ&bZ+QH\c-b.-6W_36LP_8FWUI7Z9U8AC5cR,\;QY(I1HbA
9XWSRNHZN+>8:OEaF0R(06F00MGf2[G#^4Y.8;g65c>e,->d)fX_&-)/65ROTP3b
daF42JUEUVO74G^e?.>S8@I-BK[T7K7:.YS85PB;AS-;;(T3>eP;-,P)#FSfOC+Y
/&<1B;P<C&49gd&/?>&TZ^:Mb<&b^^RN[2B<P,3He[:E&-)T3cbCBB31bg6:YY5P
VDXH<9NKXP7ggT>Nc7[YR\_FBAfHY[PQ#=eZ+Q&OH7[[d]_9I).4P1?c7(L(2dDa
#+RJV8[?65;8_7)AUVU1O08I-=]ZVe+0>-/N>LR_^CT/0F.Y2?,.X2.-d9P>+S\S
)WPM2gQa1FdBgebH_a&KM(HMX)Q@\Uc5:T_YJ[Tcd)baE^5?2VRBSP);aL[(=)C&
SCb(bA_.aZ-#Wf:+<;_<GQD0?E:U\0:/D4>+A>fgEGCHGCX5<QE)Xe?-TDKJ6/J6
4+9UJ5Lc-0;&W2RH[GB)W;fYXH\G3C+QI&.J2:?CX?^?+^Ic4_g4[FM;7,C3_T:0
XE]]9[Z-aDB:.#,QBbHN8LYcW0ZF=1D5-1<>YE4SDUFG_<-(:8T1Se9(&5Y[6,4c
+PDUE86DBH]W;e0A.9Z:_RI4gJOD5;A?+=E^:<;J>\]4cI>5/)UYVE)Of(5,O9E/
?P.U4:1NdHV2TY4WI.eMKV&02+TaH9N^IDS,AV[64#+XS1D7f8&cJJc;IT5#=;H=
1>g)J&/7+<6UCYc7_U@:PS3fW\C1.b.dC9[2?d8:1Q?R1fL88<Db/63RB?g2_#&5
^A39.cFCZQ0Z>IU+d=6+<eO(b2aZ]OXb+NI/V/X&Xd[+9c#49f^5Cb[f;HH#U\_a
H<5.e^KYZY?)d7CA^<7^@T3I4\#1[GHN(7[\13MXMB,5S?657P/H)ZbA@IeD>8I8
M>H[XM;;M&C5Q7#E<J(F=\VKU6K.)E\9=$
`endprotected
endmodule