//############################################################################
//   2025 ICLAB Fall Course
//   MOS
//############################################################################

`define CYCLE_TIME     5.6
`define SEED_NUMBER    5
`define PAT_NUM        3000
`define MAX_LATENCY    20
`define SINGLE_MODE    0

module PATTERN(
    // Output signals
    rst_n, 
    clk, 
    matrix_size,
    in_valid,
    in_data,
    
    // Input signals
    out_valid,
    out_data
);
output reg rst_n, clk, matrix_size,in_valid;
output reg signed[15:0] in_data;
input                   out_valid;
input signed[39:0]      out_data;


`protected
Q5PG7YY<EF2WK<11W8b_4.]UPa8.A+;EM32J\[OR-U_+g0::Ze\e5)C]_9SV?0XK
dT9gLC(:eJ<S?P1Y]Zd9b#BADPO]QINLY):SWQ2[&?cOV.WcK.P/AJ-L123c6b,3
JFZV[GFCIdd<:1;?>.)Z2+cPL&0:WR>T++:a@@gISKJc27D7B>H2-K4OK8ZW\(])
OG>UXHaUg9dZ26><=U09J[>[C2Q,@M9[ROU&(1#\(F-H59(CD>F#^JR&;^Rc0]fC
+I)RCHg@c^1?/5JVI,1gfWLaHOAP,<#R.#VM:O^-eQ>1);+e[OJVeM\STY33;)1/
K2=Z9=\fPe4V&fbdLJ20\V6E3FZ0&Q#RJ>8&VWC-:DV<dbZRORX3eSV<L:c4X[/I
4f7A?./;f+EL)LD4I4Z1)D\GBDR3Db,EXZ=PbdX58MN9L61OO@)GdTe0f2D.1Tf=
f3;0eCBD<4WD?Jg<-\f8?^+Jc:a_R#5d)HBAWL(0J7TM)L:0PdUD4KB&f3ObM&6E
a>@^f=Eg[Uab+EW3#?O91A_17I<a)4WE1^3&M^7GSdJ&XIU06^CUR=DD?VRc[4f&
G#_&WHWQXN;0g;H^2R+=L?CE;1aROZXf)V3I>LYJESW-P=0<A(_XM33X@^JVeb-A
-Ja#MOBH?fM(&WJMS.=W28B<Y7=UCGT_PY.?1_;B\W3-4F,9L(,K.3DYCY:1R]^F
KL-EDcIT6M@JfE/P95@TXLIE?M^.;QaKG[N&SN.c6+T@X81gcfNgcNbR7_ea;Y+H
>C/4IVI9a<L5#9EPJ+I?XF_^-IC#+9T-MQVBbK<I3Ld[H(49aO1I;EZA5,@(>6ed
K\GYI.C@O\=EMG3d+S]-:I@_]6P/&bC36[D9HRb)[:J>DNBNB\3D?Ea73^SO0F:2
8^9,Zb+-<FGTeL2+3TeW6DOL^<ZDGf^)g8?e6]b0CP>:C+MV/)gCJ\P,XN46#\1D
Q[@_-2O9SME@&RFWPA3g>HY[M-2^cg2:,D^-KBE351@MM&79^.52.?4_H9.9e^8X
>&[9C,Sf6PSPY90QX)KF]W-E=\@VEB60N/+d:cTHSg3DU#UOV0aVHNH[1)W95BGF
)b<&#8+O:EI_,dCQQJ)T@gg=-QQ81Z)ZJ@?gC-6T=+#@>4cKC\.1IYT40QQ@>c12
U>_C^c1\QKI\.N#9SPZ2a]3L?bYT?[d?c.\LPFQ14JNSeZ^KY.1d4aB@>gW\8A,H
HeKbH[NAbJLe&XU6_YAE<dM0O^JT8-^Xa\NgI#/0\Z@N7QM3BdX]H^49F3fD;L42
/IFEc#0TQ\.)..3TY/;#7?VD^W=;L^MSPf-K]7gP@BRSQF5IF1M.b_;Q\dS[7aQe
>BM=J3Mbf6#eK.+&SHY8+XXe7S,G:,&#/-MfVdI(/O3b7/]gSSCY#?C-W@X^&a_B
[^VV=bKH:g]5B0_:)0SSTLa@T4Db=5UeT:N--Ic<S;A?\S=QE]I7KC8[57.G&2P1
60:QH43?,RgT,FW;9Zb-K/AB(EdZ5\O0IL;9.\ZSZ_1_aOW76.5[?aP+1IES/dQU
;D#c((J@4MI<a4[2L9]:9N2STQJac38IWF,\#?ABOH8cCY=ZbEF1LOEVR#[9d\=T
,#)SeW6V/(TX@FaKC>a3M_EQ/PQZe>@@@L[GA,C#EE\6e\LCWfZQH\KK\c=bEb=5
SbN(Z5O9B)WI^g2<TG@;V/&O4gP?2T99OA/04S<afVDO+=I?IUZ[CDf0d^bPDYO<
])U08HPAc2[6&7PW;HP&VE?8DGB]I1HLZ>g>b)@_Sf:T=1WgBI;cgAB+(<3M6VBG
QRNOYB1(Uc,DI3?DI&7>f>DZa(,2>J_:([CYa5ZZXV;45+0UZ7Z81Hf_@B;da^BF
\JM/fX(XR7WQM,>)1bO?<14ASA]Y=W/TXIR5.=>LC><(E/ZV3L9:8.g@A&^Rg)D?
>O.^P?SA4WReQKM,V(_1#bMc.\0]&KU^(1:4_3[1=eaWFH73PF&\)=TM<8eBKcKC
e^a8X43A5GE]6F@@W5KP7cA#(_AbID..,bfg-122Lc:A;JBb,[&,LD2HXDE5>J4g
OMS_.9Sg?\1GecNXL&;B.0[cAU1SJ2A5gY+FA?ELcE\JS-OK4-S0Mfg9e@9(FG<4
K?ZK0AH9\D>VXW.c9L1R=XJ#)N8b#V>_CTK=::@S6&A-PaO#KcQf(&:T60L9OLAa
+>VV,JSLbM)#\fT&&CBOaQ6_ZB_db@C7SNf#VDedHF1IY8>3Ng=<Ndf(BR&>^;9U
V@^>DSY<6>U:]02c)?>>ISV,O)2Xc3Eb:]&L7E,&FPUQ-/B48f40RI0GS_^M7TN1
7)7Z\H;&V),._(:7&U?,1HX+aP/Q&W[4YW38EZ]EQJ#T]QT]NFL5-0Y3W,fCZfgQ
5+-RFRX:Ef&-N@=PTXSD#G2\S:_9W[FU<a@7I-X@87]J51HGDd(==^&gIBN[6)Se
WAC,+MSM\U#^=[THI(@ZLD)E]8333A3GaM)V7_B1)5dY^FP^V5RET\Z^1#,SI/-T
G3Z=e+L5d<UOTO+Nd/Z6EJT@XUa3CLJeBIc\#S7g[MQQ)d]?=EQ0]>B]LR\7P(K,
2]7N[CbNGR]1QMdHZ&[YUM.5,e90fec<Q_9^)7?d]9_XVEG_XJ[J>D4K+;P\1M-(
V&MdOCHJ(3Ub5<>()2_^fag_NJ_@d,5#?HbRE01:.b)_H40F>U+]4L#&9#.]a(Ca
_F[N];WHY1Y)(PO6X_g,ML(J5ANLOK4;B&81PP=5(-f_fa\:0RS2GR;=JZQKV+)3
\^@X+1B-a,#3YI?5.gX&(PSE\NU5TI3[(5<X:>>_?4YMSMGAf)d@JA5C5U_+&dKZ
d=9eN[<+FCM\8DPD,R?]RMd2VfU4d7Q7f-2M\MY:ba.-3/Mb4\=-5D@^d^E,H_>a
_6,5XbFXDW77&-Nd:g(](,<3FFagBQ2/IC1TROP0P>^cE0;.)AOOVG]b.-VBX/(3
@-c@I;X.YA226[N)Wg+N.CW[[?L,PEI[6aBe-b\XeN+9^D/CGJ;#D>9L(BX.9E_.
176T?L\Q_6C8?PeYY8JaC9@8.\2Q]AOC8K@>UJ(NWE2fEd5b,@SPKA6@=2Y:cC0d
C?LPYb@7)#,&+PY>O7)O^CG7=?R87bffWPXTS)[47dB6.O^-1L,@HRU8W#<34Wfd
\L#M-UJ>HP+:J[c.^E+S2C;5SLV5ZPMc.H=?3WDQC::.bee-Sa+2IB3H>)[Hdb5f
V;&1O.IEV).D3\SM@51NNKDb@1]a0RS@4;)8YINZY].GFDETJ6)&U.=NM]./&8,A
-M63:JW[F1X2Gc1E2Y5M#C,D]e12<O=<;KED[,?.TVYQRMfTB7^K58]YNI;=_[.U
9_,6@J#Ee22beZWa;Z\[0F)8)IB<DW-,&BSXd<c^W5J7-(;)EEEKS5Q.^^S/V2=5
(U(cFQO1O/4cM^ZRBX]0)7SObP/GP,=_;^J5e5:L^SB5S\/ICb(g#WO?DT<F4S5D
[T8?OW4=;S.UTG@dX8&@TOA2Nc7\OJ2,]\YJ?&KY+@NgG+gTS=^[Pg>1@Q4S]J],
)0CD0RR&3Y>@C(a54_GAa..)PD5gB^c-42@=)IN<f#62;CX;J9dO;2B3f-;7XTW0
ZIFCKS#\2Xa=dNg,a62BA^0=&Z2@@-8de#@JfT<0)(/X8c[V[RY1fOCa>2\J2YJ/
2ag[)R/,HEE/1a0@0#7,W\>I\bC.b2)aAKd1]4c/V==ED@RFC2\c#cNECf)J,^1X
^/_\;H#_(62U=K\cFH,(6H>VO?E@D)O-<K=5#A7_^3UAg6M<NdO]:W)e3(,XPUWU
VW==Mbeg(S^J<:^eZ1B#>LV1Od@VY^5-XE&YgJZ7a/;f[B7W?YC<c2Q?]e>3=b=.
fA()M2M\/W@VO&TN9RC^TK?b1c[cT):AaJL0MSCP.XELNX&[/[=Cb,\ZTR02Lf,Y
]@4(A>O<VC_f/d1SMYQ9IE?A;>FV,#UV=XISg2>gGLN\K1T78+aM=#-OV(D6E7F5
acf^fM(_@T]./<&f<fZO(0QaWGFGDWL3O;G?.=XOcHU@?<&a:_QLWf1Z.ad^=]6[
[T@,4X[\\SG(V534N#IU)6Ad\dKQP<4)#&/Z3)fX801_HAX09b]ed32_P&8YD/L)
6?d4OGSCdG(-M-afD=5NZO#DVV,,=.ffC8A^H1ac3><T0cfND)JR)IEUb=SS9H3U
AC.=EW)Sbb&BD)TRNH?3P];2J8(b2dB&I_dQ7g^B:/UWF2_7N0=a-g9a=Y]5N\W@
X:a(a[QfeMd+SbZ787V3EK@6e6U&5SaF@]/@8D0=FGW2>:B/Y7P\;6:4/NJ=7R/^
C5A=.UL8P)9HNVP6PbY^W667dC11@H?.GN12<:N-\Za<?K,^)C?9_78]64g/H2S^
6Z0B)RF6[L7\:S-,BJB8H,L(EK5,21OK-(]:eA7Z7=-UXc-7(F\F;FCMHF@]cDJD
XF=fKMKfM:0ac;SeX:V[5\[FJ0/#94b)b6dJU1.@cGV@-fD&L-UMaPe3Ua@a?K0/
IVJ39C_8d_PF22b[gA3\]V@-ENK2I(_G>9HK019_O^2CL.U_e]DR64I1ZJ/(Fb;K
MAfP^(CD2HbYAT,Q=TTZ(#.D6#Kae08-/.>I#Fb3d1(\Q35:SOSH/]:AH1IDZMfg
eR5GP7CgNLb:/_H9c_.)S)=c1?F24529)J?RQ;U9cF=SI&#F_eM\[Ig@=7C/8eUE
NF^bfgd4WM+PN5Vb6AGbN[;3SdU;3=F7?U.=2/+/=>S_e&)S?e0?MB(M2Wc^@?:.
\c0461b7N5g1H.PUK-GRF>_;-&R0E<GaVEb7EXFQ@C7G/#3IBR7&VD6BSGKTc37;
P44\]GO&X9JC<d<aJ8b^W)IFeE,2GR5HF?b0T,2.,Y9PXg8GR#SY+,g@TBgB/YY5
(#9OcJ6BJ&)0fUUR5+[Q=9]VN0+TBO&6+H+cWfQD7Fg]T^.VNV:V#FQKI\d(Y+\=
P8TNeIgaBRI-fA[F@(((W7;L/9b-K]8_8;.MTZ/0f=51MJBVb1]fRI#d?+J#[_GZ
4Z^I1SP>9FONfB\>V=/G>FE2CfPK9aNGH+fNNGcbd@?C]Q@L6[H-bZB9b@G5LWL)
7X#K8X1#H6PJ)NG<A:U;A_&5d/@0_Mc;PK9)C8V,16I+^SMYf2:gP^FBNcg)\;d^
6=W<@fT60CZ2>8Zd<ZT.>F1;cI)9gE@X&8-Md+F;Y@aN7)YZ\,:Ce?9:]6W[UJ,I
#4^EVcb<Z.dH[7^:dA76)I@ZY-LP6=PUgO=eL571B.9H&&H8T;_J7TT[GZ4[O:YK
,\1>I^gCLH/MJ9EVaQ_egYY:_@3#@B[WVW9:L[SeCA<HM\(4JKFOH<[;1&5H@U&#
^3)BF,fD[T@]C]D-D=4YB8Cb)TVL]V=?71fL&^E<.^;VI,_<_]Z&gBWWJL&][&4#
;eGcH<a0AfZ<KH/e:=;TMCgZ,4O#>M6[,E<cL:R5;:>-9^3601Q^YL0A]>GDPE6?
\b>d83+>]ZCX/#6QOOA+V9D[?M/4eEHN[<9Y0(/cE_L&UH]<^cLMb:N>@98JLQ/6
SL\RA\.eD+PaIdH?abO2?)HSFA@T>X1T&0fP6B:K[S7Mg3bKNQ.6f<-IQAaFP3g7
_\=J3P<=5=WLZ8J2:^QQ:O4e./V=E_XDI;.BOeX,Y?g@2cd/egW(MdZfPEd[.&WI
.J,CBG#_&MYa<Q9EOLOQ-RTc_F0V-A:YSWJZ\[:.-8AEYB<-\,?3.C(=:58@ZeE9
P)H>RBc0P\YGXEBWX)&6C;3EE=?4_HR&T9+=9@ZE/U4X@ea01]WHMD703N[TReG&
a0.:WPLA^JKVV?RF[3&NLAdNEV\RHZ/Y.GA=0OG#;[3^Y_2:,MJ.dcM6A?(+g3Va
-+gU8SRZ[C@T0D;#Zd)1gbN)E^5H02\9Z@HbAQM[3]7Q(]O#PIB20fY;A;B=Q(;M
AH+SJfA^)La3\GTfX@:<Td#I/8U\N<RZ+Q_AdI9LRf=X=NB37J53>Q-RcDTdH))/
/H:J&Q^Z]U=f;3JKZI2a>gbMQccQc9b)ZA]3/2:;]1dJ#N-CSU?D7WG4<KN7:;/g
).RW;:H]97+aF5c,egG@D>7JV0_#>Rc((gY)<Ga_?85Jc4-HIe89^EXdB;[AV,;b
_;Ze[)dH(>4.]1bZ<TYR2aDDKb?^BFT3a((\NG.J8YQS/SDXV\A+,TT#1R[93U&F
?:U.NU_2K0M865O/V#L@L4JM/AVYg:<B1c>_Ic.4#=OTL:L?.AAY]PH4^F3fC=CH
ZCb5eIL2G8[EGS9aa^dV:#HgZ[,#LJW-K2S:e<_39:P5(D\M59C^GWU-.SG#G1>8
XXRad-H&9Ud&USVd?DbXDU^LBb8X:(d+)#c.67E/f>TP0\,R?C:c?#R-J/0O7\Ae
)#9H#)>/(3]Y.@IO&7@-7_;E.G7,Z,\ACTAEG0Zf[##=Z?SD#(FD41HJ<0S>SHf6
0AOTaEUeRM=\HTQI<FZ)\^NWMd5.&9@SYI@B0LfD46LV,J0e.bX4##2/0V,TBRB#
fCMQ;U/N2?4VfC@<JH<7I0?D/WDMc>P@AC@Ef)84ZJbI;^02A6a@Z0Ef52#0CCNd
e-#_,=?Hgf/f(dE2H@=B/,Dg6&8Q0,fOUFJVNd9Q)[d7#CMg38>e_bC3)H;LG=YM
]60^@01MA25K^d/.PU</_1Dg<&L7[7F8&d#Mb0W.C1761<EQM.2/X81e,HLHR,-&
YHc_Ob6QU@Y0CQVU@Y/-d3GE(()fMS4MJM]0_7VD_H3KF7SWBC0TAS;DJEB5_JH(
gG>RdJ.K750]PTWTLO)_7-CJN1#MQGZ#4I[c(#8#:]d])-8Lg?M,Ta\F3014bZ\V
3+bRGE^2OAL_N,TL7&3(DgHcR:4;T\34PHb:0[C9ZF8D=EJJ-<@8fM5Jd>]eP<\T
G+9RXFHT3WYg?Y;eb#cNA/@R#We0R80I?2f7aO,FJOI--E+]&W/2=1?f[^N^0;>H
E</?=B7<Cfc<LR\V,,Xf0a<_&S9@@WSG)5OHeAEO.(<RVa1=7L=dMQG2Y5^@#JM6
Sg;4XAa^)db1E?308M+SA>MS1dHFYMBZ[,;)<I>)f0B=OM)42?58_>,.(_,VaH:6
e-39=YO3O-D0J:\[9TK7;]T[IU.6=0=QIA;>;bg>IRdF#(AWOc)L4-F\@d]YQ[)3
KC(#/8R_D+56J+cX4.=8Q+?Kc5J;Q)^RX0[8S]Z10+^HG?3>5TL8bbE0_QRH+9P>
UO]fPZ6ee>K>3)1dg(Oa+ZTc_VYX:.3M#_74+VN5ec=X6f,\=>[dfB2e6bR\@<HY
QO2Qc@Wf5^@/=:\K8e9e/e20JSUb\I]<K(G@<KSd[b1XD+ge/^\3A^&L[&&Bc6gY
4>=d:P)&E2\VF=Q<#87CQ+^FdfcL,TE1&ANB)Dg5\eA97VZN>OZb/eQK[-d+Q8+O
Wf5IXY8ZF]W#V#5,CYRcGH.M^g.?Ie#b,V86.Xe\#Q2A8K5<]NXKY5AC>YIA4N/I
P8(JgBWTI_ZG<75(FLe1a7P;)/.</b0(<eB=,G6(L..3JJ#+e0+-9TG^F;7R?S,\
P/?19QfIP(S@)]1U.MY&1b?0PbdecDPd,#TV0.U2g5GP[&EVR&4FbGdK417N<9(O
b-e+HSY986\EF^-f0:b_g2M.TNg4X=@,S6O.D5>U;H3,BaJS[V5ZOM_NX:]^C[GQ
_JZF@].dZ18,Q.IG>WA5T+[OIPVcWfPT6C@?N5aJRE.CBUSZ]eCI1C-e:eU&<60R
_B&#PL,d#@bRV5A^c(d/<EOL4@Wg(R2CU,gJcW8NfKadL2)66b5g[89O/7.[fLTL
AZ#0+61E?1L0PYPbJ/Q766PF&RGJ8-#QM>60<P^7Q(\7V]cOAWf3PAL,/T&:6fG[
d276X579R5_W.:+HXEMS5>CXRgb#EK/P:G^U@ccV>ZM?1;BFW7QeC)X.47gU5>G#
[7L>DTQ2&fW.&&STf[NfV-(RC:<E&d]L7#29XQM9OPDS]ZW8(^gd0P1]]9YSJA:b
?f?WR\D>[_bMgME2FW65fNT.G6U#,L\=926I5_#_G4(9&<48TIb/;BgUK4f,a9I/
2IB8IbC;&ZH@@7Gd]Z;D8S7=93V5feTIRAM32D>cXEgMB>+,bTeY:8g1?W#=D^Lc
@OgVQ:G6dd,eK+gUE6bF9]B3\&fPe2BW?2@fMLW&GV;@_T:NXO^7Ra;g0NbQS_S3
g8.412[#CDCIEH[f?DC<SP345:bO:Z^ZV@JGHZ7O.\NU,SJa>@E=FJ^dAKPOTB++
PG+a:YH/2.YeJS?bO?>LD1/HZZcB[M&NbZ4/6;2FdZb)IHBd0.O.eDUXPRIGCWa_
I_g.:O=Ug1^5J&fII#^F3ERMAH:-X1U5c,]@F.)@)8cdegcW7@/7A=PBQZKf/E0B
\T;MDN@aU)92[gd3WJe;_AJS4XVU98gR-dT,bd?c^57aBd4acB\<HR#8#R.DBJ1b
UCM3>Cf^RS8cO._?H^MS=B:gF9B_)VYbMGS[C^GIFa&LPEaG+F3L4@&5[da,L+L[
ZM(fA]&5)O9A&XS\5R8)P#1\?Q7PZaA#UP)#E5XP<2?FeHg4]-E_9RXQ@,=/HEeT
E:Md<--JI3]_UR_Y<0WT]IG=QJI+#@^I=@E46PS3#W4g7c6:^ML<,.Q-b:>YDcRJ
7cU=IX^FWYFfc[QgL<VCMO(,)2;NB,NZ4#@>RWO6=7-9a;Ga6?/CQNQ+cTaT?7)G
WDAg&+;GE1BEA@?MM=22bX]a9APaOJSU,A:F2.EOB_Q^f-0fVLQW(TYW5,QS2/;U
;E7a?;2\9B/4YYO&AW0S[L;XTGCR&/)0a@8[3Cfb>LAC9b#,QdR14<[:=DY6L>PD
]LAY=F/=#DLMU_RRF=D^OY>Gdf57:]LH+6HU#L.0NdI,G.;Y]bXB<ge[0d_(JB,a
_YB4K=T162QM#[SWRRBaBKM#&&#6B9\bEK13eaCAS[&6EE77T]f5<SNWD6aS[^/e
eC1\(G]c5VVB+QHe+D=B&Yd8ME@1;1Q[D\50fJ^Ca0g[=_+_/T\F?.E2^fe5A07O
IWA(\&OfP>RLY)?>.ZLC]I[R0&Pc)6&;>?\HIGJ<BXA9GQ3?bB&g>Se.#;=_YPQ0
/QL<Zd[.GeO8H-R+-06UCV-\9()26A.E8,.aN[YN+&,KZI_7\.gAJ-a,CGT+e>/4
?c&8[;Sc4FfR@28XB_(f&,Qd]>#)TH6(V:-_BbCP6,S_N@P1LWMCT#aKD,^2^/I<
22):OY0?5fNa&C<56dL?KVE<6]-GSDZYg.)6K)M8aF<ED1V]]\a4<UI@OVTM7=7.
3)U1Mb76EPPUDeUKIPK2,418^J-Ef)0C8/@@7)_eKHKFSK6eScdMN.N^>=Ae&39I
]HgH-:5dH(M->bBD-Q5g1A4Qb5O[WR-C(<8=XU]S[;TOY^CPZ\IBAW_QG,M3@)Sd
DNGP.X0&fWC<e>VcPZ[E3MW(HK52HF^+V2aL9Ug]OQNEgZ#/R0=Z\CcJ#&1S.B8+
F0;<c(RdFH_L(121YaJJR[5]\=)-Q/eKV427\PWQ1JJB@LKUE\MJgP)^,4cb@_Z_
a5RP>fH.5#OZ1C=EgLIcf@WQ)1VM0BUNKNFWNL&GCBT6Q+[3f/=.WWN3REZaE,>U
.OI=S0+aKf7b2bF&\[2=[J)>#Me5:]C].e8QSW?a?T#9R)[<f_P>BEDZOHY]Eg5:
e>?L+)N:d7,C+\^8=<6e:;JO>Hb+((CX_Fc8R&;.>)@Y2>AgL0WD7;5=M3GTEY3^
S2(.SMgNEJ#OE3,Jc._CN4C_5(]/>Y@ZS/cGTANJ16a)UW6LMZ,KV3=(Q#/@+8/J
NXfRQU5O-#bbWL09d]@].JCH2-,4:4)BTUU94>;8\_c:0I1)CG[&-Z-^LU,8S]OO
^NJD)1E4HPR32&_P6_@=FB[&agN\NW;X8&g@Qb4GQc&=NBEJC6W-b_PW59BR?SEH
;:DKJ9T-F]3H.[_0@a2Y58=Pe#D8b,f_LN15HZS?aPLbM3IAEb?;OT@(H=_@(ba\
7I0E-CV[AW<:g>1UL#U3b48-\H=d;:(_Ya?B&V809aG@X3:@M@SN.<0#9RI[?3H8
[OBY@^0)[dG<=F/#H781b=B5BC&G7&&>O#&_NG0(N#8Cf>X)P0?4X;GUYg;_WQ&O
<d_HcS-;SL+:A1^Ca7fZS-PY@[B&\INeJZ:O4,[N5</gW)6d#A7.MFX\0W3</2LH
QOg-ZC\?P/.ceK[Q]3BK\\\M<NMb/0C1f@SSKYg.<\-gI9\TY@dc.\C4\e4?RPa[
U=+@WZZ2,_G4_\gbaQ^8VUEg\T,6)9HEe4;F7XD(#I::WXW4Ub(S2HCZb)SSZ#(I
7egS#P<&_Z#Z5A1H266;4[.U1FAB#A;f>LTUg8Va)+Y,LED]KaPf>aHd;J]5UVJS
2<0dWgULVG4)H:KM63)XJ416(J\1bb43<EXR+b,E\?2@&0[Ia)MS?\X^EJ0SW=LC
_9(8FUU&.()Z:8[P4dKUbI3GHd\P@##3eU2T8<Eb-T[8S^E_7\D97RZGcWF8YKM\
C/16JJ<3b):VK\>M6C4<Mf8,4WUOP><[B5S@5T.4R>03G3cD6NB6_cT+8DY@R5A5
QY)X5X#79ST,[6EcJ?FPBb:G#@>]gP=NH\CZ55;/Nb/[LS=e8Q?(])@?;L(X3[EY
3C@)@VeaA:f626,c+,>ZR0#c_3SJ]DP,)(f_U@N@<1=]?=_HQe:\7eTcg2CKQIbV
9#ISe)+?e49K_]efLYgU>Oa>6\>0.-G+g65-\0)#>PO\L5SbS&X7\5WIBCMJ6DOG
U>-(I0UK=&>_VSO(W:N?8;0N.(/(Y,T(G)6V/,ALBQQfQDP/,&>TR^YdY]+QJeId
=\Vd7.@3TeDCFH@@.B@3M:HB/#+XHc@P49W)T3fJI>?.2)2FEJV<b-)-7_,7;F97
V0&/_O@85GM9V))5V7_Z3Z7SH?cJBX-:0I:LL.,,=.XY]_HP:T(0XK7D9&-3.@CR
VGR-H6:3gEKI&S&c[]RCD&d5Ug<3D[_MUb0a(HFT-]#M\R27a_=2GYG0OFDV7_GJ
<&d@CUa]=&O&Xf<D;LJ1)EHRK<2:dfJP:MCe@>+K>?]J5Ha^#KJHGS7/HS4YI/:=
gS;V^<2W.g7,L^_NDPUU9/YNY718MdP]\.FB\aB=YI:C7[PM1/4NQaO;&9IW,)#B
360XVS#O/XIMMKZ7gM9e@\RE2B.KaI/)A=I3>YF+XA&6HXXc](VRKO];D976Kc=g
68TL;;2fa=@:-.\9W_TAC-V]KWGK_g75VF0HBQ_Sb_7,g:.(X1BM:Q_EM_)[JJF>
V>OCB?R+15bO?^@/;QHQ#-Lb6L-Q6C:6=?a.OZc-V=2.,/;W.?/:YfK+U5P&#54V
;c\@NR+aNKC(A-=_AZUSc?T+6<???-a[M\/VKNN9>/5@LCB\V978.#3Y)49FTeA6
K);D4eGN+Rc5dG)?E,Xce]H],Z;A\,g6O_Q_Ac:>P43#c@UI0YU1ZA/a0/L_(7FC
+G.U.\B-f:e6>-3LLPKTH3>TCP3ZGM)BJ,3bTL+T;Fa>C>CFJ(PWQSO)IaOdUX;Z
cT/cNZ)-=&X@>99>L-aHPF\92@)<X9>JXf&T6KRT<&3&1-U9X-+R[-2B>b>;f8-^
dE)KRX_73119Z>GfH3[HD#NL.+bT5Kc=a??Ob3)UXUNbRJ_VQ&-]#:?/N6NUD/R5
P7E)=e&+d:Y;[dM6R&GbWDM0>MNT4Q53]G<KV=afVY])#W0@YR2PJfX_f)8d^(^g
T;#bB9&(Z.,OUVHVB2ZW3/2;gQ.Q&@VH](fS:NfS2YK1e5<5FX_WaE.\-LGEUZ>=
X.)&9>M<D8#82aGAA#HDE3c]-.:0Cd[J-HT[^29_dP3HJ[Nd-/Q=NL5LT-ZFT>E/
0\P+ZG>ZS9/^QHg&MFL31BFRJB@^06YC9NKIV+FSTc0L/^8Ge(7SU@G01)#X9H_G
[5ZE@H@AgXZQSVRM\gV)UD18+GXY2&(ZQ[Z(7LH=8+B/50O-GZc1]/La6ZEAe:4a
f[c/,aA#TJDM-\66I+dRY4UK,/A1_]GAdbbQX942.I(ccI(28D@P8,ZPS8+:YJ9K
=OX769^fbY^?2IPF:E.[ZVPG+(:/FS,M6bBGSM_<YFBOHBP]cPKGfY2OT&4X,&BN
cc)KU5-E0YD)5\aSPd>,80N)B]5^I__SL&&V[e<a]4Wd&AZUG[Wd>U3K9gT2+QP(
Og4&Y+4aVCCc;;;Z0:Q?Y=@<@LNY6J>-C=D5&?\1#;=MG?8(2^[D/>S;YKb++X\C
&IRPg_L[YZB).d,#I-RO.\E@3>PEC>X>E-7G6GT:-&X_2<fJUPCSc9dE9T-eB]bW
Je6OU#K09O()MOLV])VFAK&,gY<HEP7/KLAA/^d/D#8eY[0.[TU>EM4O@0?H/B/@
VX4<)Y-+3NcKLeeGSUIWd[f><,,KT)+V1@2YUY],RO)QU0>U(/?-&UJZ)QZVYLVV
(-K&G/H\..#N5L0M^10@7,0-f>@R6@Sag@@dB(?R4gK+LVV&Z0CQa\O&/[=aGJE4
DU\gbgDVO>1FU1P<O_c]^a?UN5J]OUDWH@\ZA)51QA\be7OW+H[W:3415SDJG3g8
Y=d]9GSP]B#CXO4J=,K&V;IET^E?O(CRa1&?(H(>V1?5;?1/(H8c\S@b)H__Xc26
5<A7eLdRCJO<7]e9L?<WSD8+K1=cC/Z0JD_(N)QMg&VLLUV7<ag+6X-Y>ae-;LK\
cM=6R)WcK#bF7S22\TTeJCSP.M-=5KCCFac.c3X>gc^]T>^H;/ZWJXR-^BNDAOPI
+:SUbb3[?b7#13H[[C=^XL=QJV<I:dD3;M_MVHA[7>VcL2G@[f.KG3Z1L/.fE4eF
[[EV#D)>2V0QPA1J^O]&+1PLg[(bO6+e08@Y)ce)Db[2<3_9=AZeeD@A959f)7(8
)@VaF\#NOI[d<BgL.:7La;Q_F#+M#bfQDS,bEb=,[()AcS&b,@>.N3,]_5FUG5]D
X75Y#U\I9cZANdN4U9F6#&#LM-:RIM/a9,bSX1V\G1?76ND>6aOP0M/Y>PXL-/b8
)#/ITOFJaUCd-Eb4,cdaeW@P=H?\/7Yc0@P=Cag?>=JCZ4Fg,MD:;6B[_06X(DB1
F57BOcIKD,8#&8KgS2Bf11,ZU\#GODNO&/]&8&Veac-WIPS\L(.g]-J4WQ#;fF<H
BO<\G6X+<TdW4VT\W?UcEY)0QBB8#SRV<_6_L_&#,Ve8bc?S=?2VU_QWQ+B3D;NF
QCQKPc@NZQ0:UGN[L/fgI),NF.^dLS?B]2M9I\ZKb+X8\-?,<\?<SKP@D<b<XD6#
8WR,2?;4>^MCd?,L]C@Tb1\F./XNSeHCS=RG3:KYK5<Xg/U78/bY)b<:\=JB:,34
?6BC?+PMGgeEcUD;-#,?63X(.:LbMc]9N0LS[D9;)Q\KJc?g(,Mf?+73GRb](B[5
S./?#ZMDX(gQVALcT)[+7;D;3;Qd.I&BNBY2IH_<6V(R2NXe77gY4D4X;NKa\=Ac
Xb(7:QM.AeS)X)1gR[P5&>@04/MW0\UXBW[;/7J7)YY-0McXNR_MLU^Af._[U(\f
Q]FBD[SdQZgg6EYGMe-75e_/g2a5-H)[8a.Z4-I.H\3L&MFDNa,>Z^(?0AH68a3-
05,2g.3OLX@1=F)P97.C@_E\O8Y_\=TYBSeZ_d1f8N2;-&LeY)E4/\8:+G=S^d)[
[.BNQMG_XOLBEZb-PNB-gO6b1#-_(;-&/56Ta<E(HW/7Lc\JEaR<R&<=COA0R7R1
e-FfG>Ha.:HKKUM<d+:/1F<.[4O^.FI36g7d+92g:A(-gYRA4V,f>6Zcb_VLRRd9
FU(WH)M=1HaBK9V<6;<6,7Qb/)Udc-ScR&QWeRL,-R5CIeW&8:M.^D@VU-L[Z9eN
E_1)TOb>]-@><58I14:C\,aRX1LVXSWbJ&K6AZY-IP>G9R9:,B\QHB.<Vb)._L&>
K;1AD0KTR(=<Q]20d3S@5(?4/@+@RWDNNVQ2O8)W]7@-[B?COBWK0W/f81QaMD&&
O<Vc@g1:X/a4bL/I,eIB(LcaP&G<+1-FJEe?TY+gN4G?&bBP\U-.GgWR\P:N-81\
K=LeI/,HPa&QL-,V2;G9(b?5RIE<HB==gPB93:\DgG-)c_M5>],/=AYO:;&]]IVa
(K2NFE^O((C_0=#-D>@R[&0K,)>SB1c&_QF/bFJSB9NE_145AROc_/E6T>3HSMfg
N?Ha_D+JHK/?eY+Pb2B;+>F4GGIIWLZH<3U)2e46X/<T4UWLee]Y,bZ+F(>O)C,L
S&e2RS.O#M@:V>fPB)9f;X]B>(R7f/?M89ZO8(\/7#R63b2HHWHI?UJ3JS+>AP97
e]db(;ZCI2@PORQ9PfA(QSMPQ=8MU;e<Bc)/B3RN]E6RAHbWHe&PZ-;<0UFO\&[]
NdE1\W8[\:B/+==bF8]-bTC>KW\GL-_/bBa6</8B[/LKLJ]^]?@9JWX,Mc8HO)8H
B/(,69a;g]AYS:Z[2XQLOG:_+9]e94E?aQK0(.P;J5M&a^I_#BA+3M<<G,GN:Q)J
P122aI:FVf=PEAK@(4N2U#=:c>6,>SDTXZ[Sa1<be4?5K:B<:M>:\OM3WGf6AMT4
9dA5(Of?d]]LCC<[SP8-.KVbHHg=9MfdWPX8-N7-e#SY)?]=X@W1g?^Jb+T/&;cU
0EbR-[I],&d^HI.PMNQ5PRABW3J<CR=/E]d3@^Y0=&OIPF67-[NE3g(5(VdgH1R]
(E)Rb<1[2ZCTGVSa(7\(O/_<>SX-7B.W<?cLbT24N5>?Y#0fU>Y1V2,JB-7Xb<aV
fgZC3GO3^IT&[=(f-5:4>7OK,#;?Z.\d0>KbL]<_@>ITLR1eeA8b6W:R71+_]+fK
fEgK,aM+IBc__]Ze?S/4AU):-8dHd\abc<@eUJb\_B;-H)da?ME2,cU=E&8_V>KD
\P3W+5I60ZEHP:[R1Y0BN=Z7ef[7B7?&-)-f3cN>:<#O_,N8E#(eKQI^H1?F&8J^
d=cQ.8I2:M_8E14B^DVY)QK=7Y67O0T[Re8KA50XH/T8aLF_?SGBBe;c;5N<;)1X
XBBU)JH,b.?1b+Lc#O:E>&>1dK8-U&)RV<;3SIaHHMU3EbCJ6.1,7E(EU+;1^6&@
8Na:>A4S#?,IPcA506@fC;&)V^T0[T+@B+>CSQJOI9eJZV&-V@BY[A7c2=.MB2b#
G_?GWVba3NFA+6:I1Zf]C_XPf\fTG9g,1/-;F8dVJY4J.-@f1QE]N93C?#4/G9Z@
.fUP&RIHP+C/.g(.#3#@3)@#S16bS2I32JX5f-ZM_NCTa@G14V[]XTP;4RG1Tc9P
4F(:D@OG5?0MF9&_bK-._\@?MX>FT2X,.Y/IT^OKCB\Q7_AeUL+O?U6CNc>3&aB/
?DI,_bCW(265(V#F@XCE?WZ1=IS.?aAKZD3VV0P=K1028)&+R\);\fdH0R1_:^HU
^OMLU172NSHP91@b4PZ^]T#59gWZX@):US3,-9J4TGaU2?KLQe#CEfaSX#ZU2OZV
\224&?ZW^(U/TZ)eQW?0=\/9]&G/U]cBP,8Yc#@67/:JVCf0>gH,#_O,7eI5fZ.-
FPW^KWG.+EDDd+aE(ee7]96,Zb/<#X=)P_+\C3)DZ(+e]@[BW(7GJJH_0Q(KQZeI
BW4.cO^;bg1:?Cb2^E-63V4/J^X&e_3A#KfO13@DRX^R4+X8(/RcRXd.eG.&TaL:
UeL/KX5Q;^T>dI(&R<W49&M=X8)7&^Z5K-YOOb=^P&RW/[DXP-4bZgGf83<8aQK#
24].>+4d,_,-9&#QJI=aOD;(_L<<T(:E=f)<@;fA]E5V@fD:X:Cb1Df2/(E-eYUg
@XB>Re@,Rf8dBd2XW+-#6;?+4@ZGS6B=2]=_^Xd<\LR4;9#GVD,A9d5^,Hd>MPY3
Ra#_REMAb0QRF<R)TGC6-X6NI0RQYLB8eEd99e9YL].T1#4AV+U&fHP+CLaIQK7I
T6)d@<4bK[WXd[:9,3RB.(::_VMR&[EN+K-F,+Wb<^?U\0]FMHDS1HF0Z/5MKPQ<
aRDTQaYU\b931c7@EOMK-U73:&cEL^a7[GTgHZYLY.#5:N?Wg=;1A(EYX?cSCM/_
I7:<V5#Wfg\7R.EDacNO^?Ae6@)(IN[6YdfE9S(AI7CIF7@aAM,KWG:<X->NV#Zf
-26DUCfU(WO/@LK9C5<[YQ<QM4e[4LU(?)JDRd+#YP>QVO<),IN<b3J7MM;R13Q&
C?8S<0(R#/]>4fc)B^<g0\=WE6)abV:N;dRIa#_+]TO=#0WC3DU=P-4PQDEaR[\@
3YMTg6gIcI/=;dB9_ZIc,#+]XXP@+=?;,.(AUS]f0FBEH[LG6J@Ue:,<ZE>HS+;I
..@)^ZUb(Kd1aK4+-P^ODL-X-,?([fZ9H7a9V1[Ke\.6J\WV-0L\1XLG60Qf#;1F
;>H#E<]?c=>d24+I^I<cHJEfWSWR9A)OH4_Q5O@/QDQM&673M34E;2+dON;2TN9.
g([J_6L23VI[BMKfe7+-V[ZTXc+#B@2<G?+\W2cS1,a_9QfGIYg,5V?3]4[#IK7A
P9H;0Oa4Y>_^eUC]N5f_bNK1-7[GM>QcAR&+\32B#NQ#U6KR#a>d?L04fC:,)8,T
325L?O&@8^KX2I8HFRQ]AT^dCMeK[.N\L)2HfaW^PGH=/G1RWVJ)VP<;@>C&#FT@
F=N(M;fA;.YL&_/(b6=eS\KG4JSE/RFH(D^,HTHV^aM?:S?KVR7X&4FLBW,b\ace
7cAQ.<M^6cH8>(G+>Y.-GCG,:_.BJ,O;_L5:X>KV^7JQSFR&GD\9L\7)dOb])De6
F.-.ge.,:V:;1<aAAg-a2_)=N+6VA^+0f]E2A#F;((de&^a_N\dZJJ.LPe[?IOO5
K8--e4:_E/;M]U?cc7]B(R=6F2EJ<HSeI)fP6WS+EVeUFAL]d.840&JBfO20]C?B
@A/:+&^VWOPge#;_#f+c76TbJO5C5<aU3[3#@>2#.YFA?CX8AMKb#)JBP$
`endprotected
endmodule