//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2025 ICLAB FALL Course
//   Lab08       : Testbench and Pattern
//   Author      : Ying-Yu (Inyi) Wang
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : v4.0
//   Note : PATTERN w/ CG (cg_en = 1)
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################



module PATTERN
`protected
W3dTRCgX7)DH4B;I>(I:F?=0e<:@#7#I\IY<ZO8>A2MDe#^7e+R4))g>6Je^V[<3
dU37Rb^UTEAPFR=T54Uc@[I]^71[Z/N+_@(?_^JE3NV;MKC77=Z#S:0fI:H2\O#R
_R^^=Mc.<W#WXC:@Vf(&>Ne]U1::K7R#&Fg#6f,.I@P,6+\-GPFAIY#gS&cUYUTM
1VQ]<95Vb2#-Q;JaSYeSJ0-O/:6#H&]Y-JQ:A.Oc6H+?c_F00AfEH3@_gP>/#9N_
.a89&?<SZMNYMT7H@#P-=Og[7[c;F7<^YU@aO(&Sf_3bGYF7AY)<0D01E\=gb^-Q
>JcE#He7[<S[#93G.Nb:QX3J]Z8B@c2LQf0c+UT-@g(X+5[ON1-1(5aE(/P[XL8,
bAXf>E2K>dcPB-AJfB<T8g(.BPa<8LI,7@B-W(+:ZODedeUYe578XMKLI0Nf<FE\
]D61_&^G3,&dG?&(,:ATJ4DZD^[gaL];W2Y.gaAHWb2S5^E?55)=AcW<cLKJE^T2
6\?.Yfb.DF=&J7L>S=42\]F]g>[R]G<EH-UG\@,cPEH5;UaS=,P9=eC.f2[-V#Y,
S3X]b>c.Y.#<IfO?QM\I5cH#WANY;@--D)(A(]PI[#.PPd,XOd@X^dfY5gfUB.OD
cB\(;J3-V3XAL?=)BGd:8#CALXP]^X1bg+<2P>M3>4CaHcf\P>Q6G@<T,R1dQ]Xf
8Od@7#Zb?GGb&gKGESbea6W4+\76B-O76M32+Z\PBJ7JAQb?ZLTWS,/>OeaJ\835
QE&>2-47I?AFRC;E-&bW4729dSQ07Z3,aYG-FM/g(HgdRg7XW5]NB(>=5a&.9:M[
U34Z^VO7;#7D2M&fZ5T8^@Ib&a8;/U,H.,cGS0&Q-e&;a54c+FJ]7^.7bOD>d1bB
Z+U@[@8BC32FIN+A4YNg35#Qd7bcFVc_AY,,U;1_B9V9GOb8Ncc&5H7_)4[g)::V
f/JZKCJFS,0NTg_09DHE>P^DG^,bXeY;AYO;A++La-gC[N4_J6DJQOVA@FIGZ,+I
U2YR12cV]#gMTR93#IBdaBHIJBJVD>]4/CFPCI(MA:c<4&(D+GSLE+;=NFN/A&F/
5[FGgMX+#F3-dDY,/ZDS>:6F20SN8[9SCLF-F_JSZb5CVc:99VWd909\N)gHU:(J
MXK?G8O8?^+U2BR2g9594gd+I0>geY+6&a>?[9-IPAc1CLMCJ/A-_T<HPME-NPb6
6Z0V9f(FYUER#(ZcPC.6bO54ea]]e52^906&&+X82,H;8KY0.-EAJ;08dCM\>COL
:W6VWC[R>B=B1I?4U5EW3P(U2dYI5:73g,a]0\gFcV\[Y6LH-Og2WAZ<cH\ACPX7
P=[bKY9Y,c(Q1([5>7YQS:WecJM3KY\5UWMd639PK<77H/(;HAJ\M2B3g@<)7Qg>
F2S24D#b@b]6U7.LLB_.[GE)YX)@?^ONO-PS]c8<FBAc\T)06-W7E?CC?_(bR\cB
D84>YXZE-5\:1?931[W1SO4ID\a)MagI_=.3V&MMM_J_]cG8;0J&3O#MgEX-YZM&
d7^ZS.?Bc0c:VD-c>9.W?#OV3.Mc?6cdV02DPK@=S^A#Yb+5[YBD]E#SHA;LW11U
),(8[MYL3JGY+(=V+@KWSag;YTMYA[C+M77ebQO6F?HVN)D=b?)YV1T2U;>dY2a9
1,,#:R@:HCAI?^W<[C/K&cL(/+B39M5BAgS.><9^RX7YA15W7NJU7#O(RdfC\PL(
APC2b_F6bRaE)0a,M@1QO4PcPaggZ354d-FZ[8eV7_FAIgY#5-?;c#b#c_+ZMAYJ
.G7\G1B-b0SRGe\#f6Y^W]PANbeOc170Z1U?\YR\S^?W=>\5LRCU1gUbWba>2TPC
QCeD^1FEC@eR@O<7SFJgaa_Y4(^dUJ^,4Qb9=Wa1;CB?GJLe#=^V#SNCV+H_7L>[
c.USDVWRH@(B10&Q<0M>;^=BSZ.8H5E(:)9([-bEgC3MU^L]AUL/N+UcB71Md28O
(a/^MU)aZV[@3OED<ZBAF(\/:E(P:OGE6U)f79QAD[-\bdXKO@dNFRf)(>=J6S+Z
8LA)1DL\G&f4@K>WgD<&HZR-4@cVP0b3W:FI06=bJ#ON[4-@HD)C.)b:7MHf&3/P
@W[@1T_:_JdH)fbA76Ag+;3CgJg8QDd,1)_6)PcW:9,DE4G)OYYeE>9A&8TSN>a#
8@.B69JOXa3)V6Tg8XD5e144(0;U^?FT7T.@Rg3#ecN?a1W64-5^;gD-4,1(L5X9
X->3C;g.F(<+B3Tce/g2IYX+7DRVHP#-WK<GQK@)]AVZ@+eS]aF:&+W22YA\UXRG
I07RI@1+D)4:2C7)4QVPS&ZKVN7-1RAH8PVLY@5XP]?P:2OI2/2=3#Tf]@?M-GN&
:FP;_4H)0:M)R,J4O@QWK?Ueg&9&+SO?X0\a\e=J-]X9dLVOGD&CXT5I^#/&&1PP
39CO)8b+1M#G01g?SV#6@3_,:PQS@V9E6/A+>-&:HE]K=;=TJA?+U\?/Wc57-/U0
CD_@5WNGIIW4QWgRd+:BCT@T&R4b3bEU2I=@6JX#cc^c&B2ES[b],4RK?1dc?9-^
Ga<?/fWPYK@N[1XY8cG<1=/Z1]^dEIHNWK[AIFU7Q;)[;9MJ^S</SY1-#geJdX@V
TTB90)_K&D-+3@Y48V(6/d]C=WMJf^=OO&L&<;cTQ#N\UQ2R1CYD&[cA)2_2E].c
&W3#\:DGFQ_50aQddg[.>?H.Vc;O;21[]0LIaNX]f.^_M:CdMM9YU7@Tf-(^J7B.
/Z^R2S2L)>M,X^0VcPP\;c>F^HDB&8f\W5aB7Y&?9;e2f_94NA.W99_QcKL=bP4P
YG7=>?8VY)/cJHB+Y_O4HH[TO]b(5#&8UCK_b?]X9b:N^WJ#bL(13-KWX__.LZRA
)D@f40RQ9A,eG\bT7MT_B)/EOE5=FX97EgRP:J_B;OJY-Sf:8#D(K5Ze@Sba#T(;
F0WgD7:0[&/(b1=;^:X@d,)W[ca]b8DMOWZ#/:0GZg=TbDNc.&)\6UMTR>c_-gSa
\>g0#5AIKgcWeSf3.]57:g-0^eX+EP).a1eZSG7[I3#8dS9eWQD,,@Y1;@03N5\U
(d-JSM/VI\-#NXd[][64I\6P6(-aZaR^E7d,W2TZ19KUQ),DIF[/YZ]1dI/aH&V4
-LJB+cGY]X,GVOa]PTW)@5JT9AOK)@D:0WVHT&fDI--V?\O,K]46[SWG)HJ9<KX.
S9YL<dCUe5=BV&U;ebU[=A[)G^Nc.BM3PZTP/&48(&@PHA2E<#M,eRQDAZQ,A,)3
>W.O\]cYBU/0(fV9UT>E?;WIE0W9[&ga7NCad,Eb<<DE?eB,=2+3D=FUUPdTQJTN
3cUL+7;G==<VO/TdY<(]SUMe..3aH/;e.IE;LHKfc_+-4]^QIE(S0#BCK__^TVX2
?;(]ED9G&O5W,B.b[&D-T62<2aDg.\47EM.^eDV?]K=VQVD,<dE+,S&V=gX#N9Cd
Q?Y:F0QMAaK&K.,GbE^2AXIH)>-=c-I/eUGeI0P;fV&81T/DD3A:SA-c913NA+)&
)G0X9]1g\O,GM1F9E?3gCU5.E.7WSe9K,9DV<8C^BJ9CgY,H:/>8IYKKa:9JS0_+
[f5e_EgAXJd)a/>DL:Je(&7X(#b,+Y?TQ[JQGX&9<<.3d:>Da6WE_:6#[D^DO].S
=F@e0fUSON#RY)fQ0QL@]aA)VgH6YZfH1FM)2?2VN0V/N_@P6JL9#0]BCBU/>eTF
g;a4bEKW:M-(L7+@7^XG=8=BPCK\R<dNJd?,PQHF^de[PQc[YN^(+NX9@^+JO:?.
7Z=Mef0HD[]-@XOeRN_P/K.SFZ5F?Z\:]GK;g5)1R8DYbVV<8\PC,,=(9EOW-F(1
N)Dg)YTaCWb@U_C6)Z9KgY#Pe=fecC1KW?(TE0V:K[?@S]QV\=Ud_K]\gLEEeIFP
E9,7(6JN2\#(AGf^9PS.JR+Sed\.;Z(aR=eU6aL#+#FN0Lf2BgW<7A)43=gQT>8,
;L0G_N@FW:Pa&1=6cPAZBLT\f)Q2Se<B^7g>?0f2A-[bA#8(cT-V<^>7KDU:R0KK
O_2X:1-0GJ<8cGJQT]AbR8@>&TCM5]DZP=/;>31:)R1PM.OI8)EX[CH>.I^UP<?Z
]V2^YDCdNY/E<Y4AKG\7<=)17(KR1BOY^F65d8[gH+^a=LOCJNNN1^6HeM)9>aIJ
8OJ-I-cGG/fLbK#]M_3NZLP_g+Ne4O6@[WBM1VPZ7XM&/E+QHIN[=>gU0H+X7M\D
8UM4NN<dSBcRNK&<D[UHNTa87YIOR&S##2+ON;bU:1gIMC7A;IfAE&V[STgJ3E3E
1T]OC#Y+PCMMbfJC^:2(I70W=R:RX+OCB)H^Ff,^3)cY5Z;R4?5V/;B9;ZYXA353
d=M/QF513HCGF9]FNf)6@aL]CTS^\Q))b[SWGJXF;VIE^Ce>70BDc>Fb>M]WTNf[
P^TEUH-..3P^_VBMW7:V9MVB]0=fQPcc[=R;V0<a,-X6^-VeX;X-KD>_2aV8-.>0
87T)XWJS>#A\WMATJ+)fSf.CZ;,YH\M08J27X\2TNJ^&UAJ]E)f6f@/g+6K4@KX=
g()0NFeW8Yf\WVCY1BLD6Z>SOG-d?cgAbcB88.CFZVJe0fUaDH1d#fQZ:N+g98>^
Hc-SQfCNdM9LPb-\(:.Mf#C)#c\;Y0.MU#+B64TMZ,HKFY:bI4NUC0M9;d;+gf6[
8DQ;Y<\^?O?SBBUHZ8DL1ZB>>[Z9RR8UN]8E4b,dZe7;8c3[O/b]O^9Z7SB,?#OF
2/1.#IC<::DRTMTfdV,H;X3A[6+N1FOUM9L35?FWY?b#_gf=8/;:ZWS-\T[EPXT7
1HF(-X+LScMPbQ18XSHG2f>86YE6[2?fZ=]S^6@ECKRSb\>J29gg+[W/3G./2GY\
-8(_EgfU9A-SKO[#13<8D#c<P8@HOf[G9e>O#DA_[GX#^_HYXS_@DOR&DY-U1FR,
+Q\SNFCC(H4/=YWB(XR-Y,ZLLc];(XK>=R<bC31.YZg:/fN.)M4GLR^C)FMe^WYb
d5YA+<0b+\+#4AEDH-@/a)D,,VM#-I@J^=U4Ube4)UeMY_H)XW;&MGS#5@&Vd__-
X;8g-H7N7L)X<DY1/JTZG8<I\FT^@(c@D3f[T,b:0=Sg:MN06W&U&&\<N.AgVfeQ
62,c02CDVgRP>/PR@M7GWV^W;05Y>@a?ATSR:S:@a5#7M@UE#VaZN=4..DeA1#&\
5/0KL91OM84Q@VgSbRL\-:.W+BDH5#1Df4<1ORC)R6P/TX]GQ@Z=EbXZ2E)/HZJ^
g1?ZVT5-3<GF-]R;7C9D>R1VA/-)/;9\ZY:.c#aZDReRU(@11KJ=-S)5F1:\J63T
U^B:b.UD]#S&1&718_L__/K@;(cIFG?KOR0RF25F6O;,H&N0(^eg6baLEcg0O(+J
<Y]R=]gMOcdJ(0]:U\.--@TDc6b@O9c+<JBJ]f+3RN79X+/GBYR]FCJNE)QZ,Mc-
I2F<G#>bfVg;D;6]<583(UT\A/NcU;2OG#QUR:9\2dF/09]+(WfGWNK-AI+7Ab.P
&+9M?4#U;N+83c07R]\]+@]&WK)[2ZL##+I;2e:J0gXT#^]OARYeJIT]>6Y,[FcL
[a8O<JLPU;[XJ0-_42dM;:R>60X9CS9bH44(a13X;:--I17e6K/+Ae2R]aAZ9\72
+(8&[;-/(OcWO@a&Kg^9^]>b)gW:5:>EH3@\BE__L8NLFPS(=#;dSade-c>Bf7[2
632F)=V&@^2A=a>PCO0-G]g9WeQ(_5TP8F;g>[M)<I)ef]200;gD[WIW_g1FT:<H
,6S)1-FOW,[@&L=UcEES@OfHe=M<E;[Uc:;?B[^[;^cEGUA.&UHES]7>IVNd<S5M
d,#)&5E>Q3BDK);#]G[MLUC-M6]H:Mc@ZGSRbW^&BVf/6-T>JI,C6ZXa?V>?Y,J<
HY@[V35Bdg([05KTg+a)4QA7:-UB8(/b\M6Z9,aY?K^aGH&aW,A2<F[e+>VA=76c
XIYSRQf@MK+cA32/7SQ+\T;1E.EGONUC_.0]..\_8>6OE?].VG\C>SMT8,_;B&[]
[S(<C0eO-/=<Z)8cR>.OPd=X8>-/U4530)a(/L&AFG(4f5MPN3EBI,dK-bCXfdC.
aV:SQgOFB_D5\b@42,F?6[dB#P:&1?KSZNMTf>I3C_F<,@1=2BN9VFHafc/W7feD
><#=@TK:]eROXSDC-X7:P<;Y2L1N\RQG9]IS8dA>([WgaKA#\Uc?:6W]C@M(/-XS
fV?d#B.JFeNa#HMO-2dH3_Z&KJU71-_c=V>M^JcQHK@FM@:O-,aNZ[6W8[#32][)
1#,bK+0XVZ;W4,GXWDBaA+Y2B</,FG_a^3]>)I>2?8gcf>3.\ESPHY#V.OPQT^XW
H>>bPT/=Gd?=V)&52KN\R8=PEE<cQ;ICbP</.:ZE#\_&]Id)[UbE9VG<ZYReP_0M
VDKGOAa01<+:KeHOJCf:K,UV&24VZ?D]30d>3Tf6F26X/_WNR8&GJ?1#5@#8R4bM
FHbb0_P8@Nd+0^69BR](4HUDd(:4.6-_(<AU,<Fd76M-H6/b[A(;1N);;2WMQSgX
H1I7XJfU6.BU@]_GG#[.1c<-C.I>,#Z?eLUW<DY:Fac([8@Cfa.WF#@B<Kb1;K02
<aRQRaeJ-LYd;6G>Q2c_/VeCEH./U\2#HZc6S;?eFf\d9&BBY_>/I0eP=Q/D#a[;
&2_f?gY]+EYW2Z);9eAbRX^<(SRJ?X(ZVS<S/3d:LZ#;8gC;fA^H4AbI-=R\^A_U
</a>g/f9WPOMK-<G=2(HURSZ17#1.QL.]2>f0=Q]@83:K/KD8&[L@YH>Y]ZA<8#_
T:#5YT_VZ:1^@<YPb:73;69VKdKIYNHfBJDZ[KT3Y_1X&Y)8:[f<QK4C:9@.2&Cc
fFF.F6-0JQN;@:+9)G;)/P?1\/aQ\XBK4d]1P^@:gWfX\aMCH:4,b9@gCaV>1>c0
EYfd6EDa6SE^W/;52]]W12@U++^U=BNWD60fTK5a,8@,IdK0Q/L(162CWEd_CDJB
CR.SSMLXV#^2PGgSM2_&dU=^gbBDCVe<,\DTd]WKCC&UE4dXSS+,FYD:93U=L6[8
:+<.Y]NALT@&PN_#eP/;aPZH)GM)#P34U9M9>>UR3PWA>eMe_OPY2^8T;+f8B>O]
I]V6O+,B)(6(5f?AdXNXZ^ac<()DEdJW:X<Ib=YL+IEJPOc(&K\&?)D5VB-)/#X+
,_2)J?C9:Ig_]IE.N,1I5&=a,IMTDV=L_SHBM?8)HT<OI1\P(_HAa4UPeDK8J]>Y
>).>e?RS\1G:Wd2\;]QGU,AYCI.H^?6G=e9@/A0I6/&GHF63Dg44/G=U9,0g/I(g
9.6339:#L6ME(DBcLJ);g=3N9@RA)K>>K;?QQ0ge019(XCMZSMgSBJG+.&Q:<-5[
PD9e&9fENeQ.W@,TX9V)RaXOK,@4b/7V_8JJKRe>5U&F8T2=Ya>&dF[1AU_IXbMQ
FT>b6S(=[1A5M<4eg-](EGVUE:?6Fg4OR1MI#YZ.3<1^H;GNI82?/gJ/W1)\41@[
MB.L57Y4]Rb.S1a-;@:?DO(YYfA4Fb5?6EAH@I.0SX)AN\G-e)H\N<:AZ(Ib0Rc=
F?eX61[B-1,eGg9I+P.d<@2RP7DKQe3[^g=/<g<N,DDGa6A]cAc]33[EP>(#Ma:=
[U+42/J;?PIP;3D6WK1B5[1T0.G_gLHa@7/@@dYWF<Y=\QA9,^P[fTE?M@82#D/8
M;IATK?73TS>E5&YX3)<eL3_G(0[gVI+f9\5VS@G<^./[:5H5K7OaLQ#+_QP56+=
c6OdP>F20SQ45<TLA[G.>0aG.-R4(^&O[45eOP3W[=8]AB.]F@8+[:82S9_Ie@D2
.JJHD;DD=VeL>NJ:aJF1<4VP0E1QgHLZC?d\1C7#+A6RA5^GPFdRKG6=11b)RZ8)
1a55>-)AfJM>R(8UKOS+X3#U_T>G6.aZ#;L_9=Fb+867@PI4DD&R8S)(#ObE8^:K
9[KFBY+N7=/Mg,VDdLf]0;+@I]X?Q_OQ3#E3>;Y3D&3bFWF@AN<g75_234KERZN,
VIg^AR33=(=7,#@d>]RHQZBI=)+,:S\N\PX^A>O=XC3MY\^TV8RA6FH8;Tc:VK61
FAUdH=&&R^-I\,7JF2WNgN=9SMEOTV82:S79T/E4<GbC[6.I2,9d?5@FMADW3KLQ
.HL.gB3GU^\0g,EG^JMf1M1().fI,cg?/Z19/7&X3eQ[-Gf>9V(.f\A=H[6\_YH<
9+.LX5cQc4S@c:T#geX?>N.9SeP];V[Y]/)\T3#B_=G?=A:7:SD2]V#9Y9D(8-MG
Q@,Z_4MWQ01,A^AaA]5<VE(-bDS;,K+V??99;)5Lc3J7ZAB#E?#[=C<;BV[U7gDa
Ra=gUe9D>Q]B,Q0>2]]a+FQK(&HZM1A5]AfXXPSEHSf@W+@^D&;U5;N6[MQMCM7X
T<F@bNA1UdYK<(,g=<&(6?eB0KT3M&8A@>8PFe&,&6D/HB/]>H3]d<DPcF<Cg5-=
CO,,aD6V1O&EfFR97T-fI5C:5(IKZ3WE()(0]ZP5JS+)Reg):ZN<<YIAHLHCC9d@
</UQPbWS[@2a[N)??gGW_3\f-FOdW654[KNE(E_b&W=P&eFQ>+0OMb94Pb/M5eC=
_@8=_)O5APOZ7310fK7E=F&Gb>eEZ\;=B)ePL8;/M(_-V;:U:ON#:\90Z1VU6RJM
8T3e77]5J7P1X;:.,^+/_Qa9]5IAA?S]N6+SH/#T\eRb=,=QJ/W+X.&561ENd9.@
Fg_-)OM&c@4)D/c?)=72TNCbVQA6-D=:E5:F)=T.DbI45\E<>Y<)d4Z;OBQP1+JO
S??eWAeb9IV7:VR-NDOEaASH?RT56.(TG[[RN3;?V:/6=H2[R(cZd=SbDATNcPE=
#@@;F0]Nd.Y?CAB,MdbG3aR#.19.0B2U:)MD/G=cBe[e8+;/bB:&X5TDS+9Q?]L=
7S-BEYEcSW2:>XT8a[FTP;>)L2cWV)06^^[>Kd<I08[<D+a88;\a[-6<T]ND764d
#[B]eH(]^CAI,Qg\&N[5TR)_BE:DP+.#6C1ZP8&_#/7g3g06=BZO-_<)<A)Y(6R;
>?D[BF,Ha950c.Z(^B290=]_.S(-/3YXO>W&gC:#60U>=b;49a4G](/-ba9QS5JP
>(J9,#TaMT?SG<QF@0C;ZJUc3_KK=HLECFLA9LXU?_3TRYf\&:\?>bV+@c)H3@)(
-e/&ZfAA;HQP1U_BeM&6S/PR4MU+F_^,Z6NEH0a1W[9J5Bb2:TO1]gDA4S4JdP^b
(<2HKVg\HFU68ceH--C]+F^6U<-T)BR?KJUTM]4bMGKLa5+V.DH7#@X&B9]Vb:YK
AaJg;96>NVH]IgDBR8DJf)_59Z>4Tb6.9N?379VW46ee#:f.NCLb^:b+OER8=,8a
gG[YQ4/<f5U12>UK(2//-ge;_N>]_N]_GT2:7BUDC(ZR(\Y)7_,\9?d[Ib?VZ1bU
C[_>ZE7Y[)6;_CRaPGPP&ZbV<^[:XD-=J9aZL4(@(dK;,:Ma;]Z:B(UZQ3SC23DW
UDcJ\VfgAA<==f;0,e&?)HUD&LDLd=J.KAT8b_97;A9\<P[c+G507CcdEZJ:7]MI
Ua_0Md31W=L5D>MQOM,,a5f1Q9Ac>/e#2Y9M)K^]&N_T-#7SD@IH6-0?(U#>R8UC
S(>0-@S2;9HS2Y9EGY7XVC^@@U3>,P:1d)g\<W7BgWG5MXM)@dT]WG78R-c,X&;P
KB)AL[4PR2XVNGa8[8c>HEVK<5<VI1-Ba.-TTK&,2gbCS3[U=;\-0:K0IY?IAH2/
LV?@XHL-=_5UR?OU9UARf@B/]8]Ec=R6P0:/>9_X1Jg/9edYe[bWJE,=4_P_&WHX
0]20.e6ZD47g/9e.Y8]S.UK+5)JG^\\90\N:>7B#(WAQ@.I<\N66FIaKAE7])<(C
@0Y85I3>Ig?8XSDK/D&7YcC.?Y^7KfQI2P@/XN&Q[]?UXOe#2/IZI:.7GJT@1L99
SBYC[]]1Q,?/+Q]N5Hb,HO(e+R>?S>)H0GYZTc3\&I[@EJ34^(J?C_<)+Ne]R-@3
3ON-DYaRM0OLG4.J;P_7[+-[:5a>)Hg/JW=5gDPS)0G_b(gV95Ud0a+9[[D>a(_;
HT/;#:3Z(;FNf-DF;+-2#/+#PL#.P]Hb4eY<[TK^T87<^gS.ae]._XEZ/?,MJf.T
OYZ&0>M#=FH-AP0f-22@40d_HUHQ.FQ1=C1bXXbT6agD;6^Fee241<R7V18dB_4g
\[ZPc_5)^3E_=)Q[<;3AdVa@#aKG4A2OOTF1Bc^#Ia.GCP0A;4RC:C,7Bb5\PC,-
QR(=&5O/@R/:L78SB,>\5YYCg0GG/VF4]=NJVNH]SJCC0+-?fB>MQ@bIYdcFgace
9#U9:UREH^8,d0JT(YYAC1SSM[[4b-1:W1d^g]bYU[^Q^HG=,V?8LSY\^V6_D5UT
6KLV@5gXP\DWQ(SgId:9:Z4NR?=_#M.AJ/>IX;fV@P-/.)(a><f\<BcH0C\FB]JD
e.F_XR.71A]1&C9a2Z)\4#HX-eV@Q9.=BMa]M(GQ+CUT(PU2\3>J#f7,O>/7XL?D
,dT-798/9;6;?Ef?.\NXceKMO4WM/2T+W1aB&aHSB\/DJgI76+<+&WOQPP^>KL]d
=EQK>LGbFLd+1.1KZ-4\X6<F;</B6JJ/Gb4,#M-][[[b;a1^5MUT_PcC??.PH(H:
RH=TAEGdS>9,Y4J=F4V;J/=PTVCXddf1M;?CH3N3TY4+1,Kf]0P4K,LeJ1?0&@V,
M5&:?gJfL;;Mf,)A5SP:((+[g-<4LQd8e(N,MbC)a,RF<IL(gU:<_KMT&a@GI9>8
T.17;8V/K4NARRQ#&[3\T==XB(a5L,CYc,N<2F&+g,_HY2E@;3b)MaA(UW:V(Ygf
=3/5OJRYB0#^)(71D[[+_T#?f28F.8aC4X(POS-:e\1_R1M=c^IR/f[=^SYW7-<B
&P+QQ[ME9ZFaRDZV3RI82=.f<P4gU-3<eKFVT#HG++\_G3.ff?05.3R-VKKMOTTK
BZJRb=HL#bQ^\5[d]53:6U^:4MV?,>cKdOSe=gPbU/PT\J(K&<B/fO4DE)AJJ@?+
M19K,-VI<TV5Q8?f8;Ec-;)VH(gK.EHeX_7R,cgG#K)=42N6[)K,QS92W]4&X?AH
B4]69f2R0MSc6WQU&_aPWUZ&FT++?HWDF<U\L_7:d<L1Y8&Pg@:N2O.\>\[QVP<\
W+7Q8?=T]55D1Z7?^4-+)Q?=5I]:V9\PP8VOX_Hb/#c4dI&f?.S/9efLR6)_CSM^
-/R:N&RMW-#(YagJgW,H#<c2GHGNVDK62>@=4ZEfX[LYc917U5VP/gH+dDP]VfcU
WXFEedG].GML_P.KL:dI1&[16c8NeV81_8P)G26(\+]X,bTe\B09_04MWEXM,FKd
,@ULN6M2@J:a:BTC-CTJ;,S_:#bTA[]OU:]E^AJCa9.Ze3PBQeZdM)F+:WNK<gA@
5[Z,VbN,LPAYP2[=BfA4g4E(\G9?V.GdKRV70^]YTOO6?W:P>CZ.NU3aa#+ce52;
[&:JVO1L9C5YP=)b?APE?=J#19CXH_QX#V@UF7Va.UY>ca<b&YZK;bS@:6&3I7C<
2bE<5E)\/b8fS#cQP+DTOObX)b_^7<_:4ZbA+0N[(:dAL]J4_._a/)^f>BC4/aaK
RW0?G<>L6<DYQ93TdQB^=^L3I=-4FI>=HKdaSR]0/WPDC26MgN7\>_C+?e.82]I5
6V\f@7MB0(9ESP;H(aF<+2X>)9\4(VbR&gdSQ\(&+/PJac:F4B;9,ODJ9B>FKD\b
bd2b,88+PQUW=>YSEO@&5P>.=9/WIL3BCIbgcX9;?02:-X-L(#&Qd_3#3;f&^Ec7
_][RbYHc_;c9Y0H&+aDBW7,T)V1gL/5Ag)YS4aB\=eQ;@_e?e3>c7A=#EL)I(f.9
GE[\&8PIFZVGgT15S,P:OIMH7K7DAZ3a5SDQE@,1\a.LQ2=]M&;9[K[?Q=.6dDL1
[bZ(QTOEJ-X,]Jf11D,4XO+M<XKaMM,3HT<97WTFg+:6#<\YVD6<X_bg5d<aMD/]
gcE[Z\/6b2E@CX&-K.[#UHe5+FT5V/S@[:]JZf?00,)H60WgE)GDe</F]+7?3W:0
?Nc+FcE+Q?[c[)8.5e]_J(0K.<+74=JQM\J_QE.8&/[d#4LS)I&2XZ3Ld@4SPX2B
_cQL].FO]@/E>X[YC^=P.@KM#PV(\R#W8CS<M@6bH@&#HWHC9@ZML,+f&5@G3O7-
OdS+^FP>b4D7VVKVcWEIZD?Y7A.d-QU__9=CWCAJI?N4&R7U:;/fZK7?c-7/+4gG
CW9T=S6;LD@<;#MB4#),(4)?<@8g,Z(=++/;\B=_USW-NN7T+H[[GN72AZNaL:b)
OX,:)L[aV.SHKId@W]\RVDG/c&NMX<8F229<(GN_7HOaD\4:ZP9O._@HXJFY[G3;
.RdX\=bg[47g;TJ/O6=5]KTRNY(-P04_JO>+0696;W6A3c3;I_V5Y0fU>A/<I8_M
ZK;,EcFQ&5KeYX\9Z(6?47B4C\VL36RZJ:^&=L2g>&=-3N#CeL]?P^9.b_@?+-?U
#MLGB&@^NUO0N4MTE^7Y)S]BIU(/CI)BW,WLW\4PdT#68b>f/^ITANRN9231BT#V
^Pf-<\SS;CgZFQPS#a7M8&\NI<Yb8)5>[dJE@@a3V4c[dK8\gJf)[\6?3Tb^gPL2
e:#bM3[W013-6-CcCa;^cfERf)1f;a-c8IF]]PNRU;:dZ60@g@<7AVdZTXa3HL4D
[gfF/H-,dg.GK25Q69JADH5FMJd=[+;9bLfW:bRZNb.QF1G@f6g99^OY_aD;3K9N
eI7O+eH&ZcNbA<H\JZ;)#D0BK@:;JJD5S2N7YbPM/EOUb1HfgL>4R8^7I@)9HDf-
fX,]2LPfZ1+7TeUXgMM#_H@QPWK9fKfc=)1>4Y1UZEZLf[M=U_^d&W633L:H1PQ[
6?QTO10[J7SHAd8FdPB?#bB.#dIL[?&^7-R?&/9\K4<;[8]\d-^4@A\D)800f)V4
:e8<N&F=RBKRD()KMUZY0B)38c,fP0H-TK1YW?5fg1g9-g2fMd<(3bd=XgF9OU:W
4#([?URLccZ&<Q9=6LeDO)(L-9QbCN>c8\7GRNFL2=@;b_\-+5ID[W(Z.,Zd0b_X
I<F;WcEF?TZAg8W)K->5>_(9;VF<cI0G<4,g4147;b#\A:IL4b^1>Y2183&S)8,b
;3QKS)b,>aVFXMN=8#^5OddVbXQabZT6T@M\RI5d6K]TMaN/M\Le3C7KA)T3[Z.N
I9I>7]aES)aXb^XU@QMg#VK/WDCI+a[PZGY)HZP&]Ga/#.?cW6I^6<4]IBNXK]6f
YR?c/O4bSXCBOBO.PWY]3<d-QH(OT4c/@\A61M[?C29>[M&>XXL7-W5WA@SHf\bO
@@b173P5<#@,HRV.7/?YM:MEeUDg;460R:R830,Z;GGc,]EeAF_BVf-&_HbV<III
.?dXAE:3C@5_RK_CbL/]CeaDKP[:](KKT2TWIOL9V]ZS2TA_eQ(:MYNBd@=PRgYd
?A_a.;:7;\=MWfA3Q6-5(5dUEI.fH:5La10<EeLZ-/ZGdFT7a94H+.,D4eAAQ3/]
@dZXg,KN<@1E@/Q-DP.>g_B?FKCLJWBE6IKXaeId/ZNU#RKI6==6HWP;1@<05L[F
\1)^:NR.2];2Q9QFc4?ZY2A1A&V&AEg)CW1IL33_S_AUB[[4T>8:BR8<+H5-<G\S
1#_g#VgX_c_G&D]Z06IBfc-H^4-=ZM0AODY<)a?V,OD:E=VS_?^L;H0^GJHK[5ZG
]H,@ZeZUANMX:B)GTLSZ\\@aNg/U_.GJ3FF01YE+<[.c=MT+a9.=)MEIWB(dQ/UW
TL33M4P9Mf:[&F9CNCTeb/<D8:)LR22.#>#?dRFW8UaK#b0ZEbdc]Z.SF-7GE2K+
\90X\35(aU_A<(;HdA]B1e9@<3])09^0f6&Y-Fg0ZM>);09U7eXQ)885F@F^g0a:
:&;FHfg>VZMIE1F<B#>/KAO_Ad._()28GebQLX-+\4[G+EU@JTg]=;#XF=KE.X1J
We7/[f;I4)Y[-1+/>cA,HCD/NdN1/(_7[D]f?0=9KJ-W-]-P\T6VY>R^>FF5Mf#4
B+2\NL8C6R<#C8A@\4^4e4QI6RgU-HZ,aP^HeQeJCVWAag\b0/B2>QN)JSY/SXL4
c6ag[TBC,=K1JL&UGL[2g]6W=HKF<JPPR-EU.JWF=<Zg0.G9<87QO#BNVd&gG1#C
#B87cL;cB]NVHI<LcY^fC@J_//U8K&)J<Z._CA02H)Af5a;dfA/SP@b+@R.Z555.
X8W_D\dQA)B>NCFT#3(B+HfDGFF,#9]:-]5+PG)R\V[QN?.7L^8ZGgXEbbfT)S23
g6(^C-]-#a9=F]LJU\&U]()04d9<DL+@G047a0\B?HF:&Gc<&X^F_&.QW+3R1b[X
a>ORKd4,d&=Ie_AOK^:[eQLa:a;J9NeR@R=]CbE0f0MbC0>BS7d]BY&MHXJUP3]<
2aO^ZR(WFWgG9d;ZAgF7U@-^@9-E+(c>b,fd<-b\8+H(He]bL=0TUgU)Y@.=#1G#
3&b3BC0,;=IL<gB=6(D,RWT/K:G^cfR\JJYZB29NBVXM.eeJEMDP++<daL/4Ma8[
T3YV#@eD/R3Ja)ER_gcM6T-T,-/U\fNKDd0+JJ0,=3e,gf(#P51FG)K_T98N^C5f
Xf&e41]7G^0?/>WEA82/_#:K())JS?MO/;2e,W80VFL=Z40]a]F0)cW/F?g#HgQK
(]_@S5aU<a167>7aMRIb_+bA-HCMDgF)eX)BHP1Y(LgZ7ROE8H[)HWa0c<a,Y=T\
cP@73T,d2&LF,7>V_[b3-&(7/9#FY>@a@GG1L@.V>MM=(PB(JP;K2..Y:]T.QXg\
/I>Q)g\CV8B@P_-P)-D,.aLU,\3+4[1Z7]F+L?;01(J3TIIT7Tb_9gW<T<LfI8:f
#UOg<-Q^#3-:.)HY5O\]Cg>c.a^c326IM=?:L4SU+QK\MFJg)WdT^4Zfgd,<#L)g
TI\2.Y0RTUfT7HdW[KT,O@XbZCZMXM[7F6OY65Hab.)<F.)UdJE3)[&bW\+RYO3^
WG4,/WZN8@@_><G?A#S+?(<?29^N6NS&]YF68>c:/^9M\RG1^eFNO=0191_:3:=Y
Z>N6a\HSF.:?Zc9PYH7X]:RKDU,W\2KaMCVTfdKRTMD.JO(J><Ja/LDQ0)O@AY4P
Z:S-HO70Z_^\=2I6FV&9X:b(64NHD7SB>G[,&>;K?L7fDMAI^VOS50U#?,Se/O(e
B+DVcKX?..&]Z.)A\TTd(4?7\;QJ^7f8DC(9X6R/M/0-]3QE12Kg1\.ee7O[7[)V
(E#M:_/79MUE/=)PKI/Oe1)TcFJ=0Tg;d?5I.N=?.V(H\>A:+JZ/8=J[>=U.:4Rg
./c.\BO0/H3fOSe1f<,bZ7Q<UL/+bQbBWRD0.6e1VJ-fPf&[Z726=cC)+H@<-H-[
FH)R;[6M#C-3d(@R9;,dBZ5G4.ROAQ+I8-Y9\:>aEFUF7X5UCVWXW/O.AW3/dT9C
??.)</&4bcXRe#a)e&V,I3\[@F)O#,&F<I)\F;2aZ7\5TUcO1CUKQ>@d-(c0V/V0
IT8O=bMff(g+AALBX&FO<:P;60(3@_0R4[fD:dHU;3DKXU+c@c];1?;P>4\8,:JJ
a2/U4fI++>d>FO#:2P,?J1#+3,:]5I]69Z/?)_N8GI,X0D<4S\B^R.:>VOZ0=-e=
+3(e#;a)Q5NPM9S_K2T86.U<cd3(1=@-=_0-Ad1_I5G[1,/.?1c/Lc>9<T.:1\,1
Z_QAgA&[P@,_K)=+0A,I^8ETW2gT1PeU.eZE?Xga]\dVJaAV(\_2H1Rb5;8/XdSV
MS9I074<R/Ib=Pb4M]/D/AfgX4aH&5e#)6=ZS3+Y11;CB=/(WB6SSC2NcbPPg1[0
H#62D-.b5/Qf?<Z6DEVX3_\:DE[BBPKFV80UJ8S9G6AIXJD6c>RN8Faa6f_CWF3I
PQ:-+_XJJ6(R7UTaW7-F\SK<f&dbV\@B1:M=8J(ReB2@<eC&SGR;N:c#R_(KW.g+
NWMG&@?c&Y+.L-QT[KAFOE<f74XgDL7#DNab8<&1XMS-69J^2)aJcZ-L)3MPI,JH
XDYe&\_E:CXZ5/Na=H(+C\]^e9W(V8BP;]/:FcR58.<:NT-g@R;bU/9PEN(;P&=c
f?K0MfgN69<1F3_OS]=Za_&f+&-NY[@<QL)Z.7Wgfe9M#=b#??Y50_2M/[Y-bS]F
C<R1ZY2C08EOB;=IbNN=;4VfYAE(;X^;:;,=PKd.)-@FJNRK>OLO/Q(4bIE#-BF&
I8L39fG&e)/<RY>>cYNEZOC)XI^Zd.]b]Bc>fJVKaUE.=Sfg3E3DMNZW@aS57^eR
O)SF]O]XVdbYf5V3NU;R5.U>(R3+cX]YP42YLD1UX)Na:PgdeC4Md<#[/YO8(]SQ
RN&7]5V8[_FCCf;KbJ1)915UUg,gYM3(N8edccf:4@FGD:B_:9NJ5cIBS<#JUCg3
5GAYX0H??HfK84LZX-GH[B6EC7V16,FE^167a&@29g\;gDJJ:/QdQ=H?WL<P/WNe
_H1-2QG&e@=;9Y\fGO5,Z8/^@P/G(UMTHWXN3+b2J7-^#F.b[8A57^KS:DVS)VU+
FTJAGHR2cAe9JE.3;R/N8J-7&U(K+]g?5M4,MK@ER\;>\+>91<=UH7TeXd<K5<JN
)Oe5WBW4^2Q8^>62<CQH<+aUJ[ND-\FWc;5&R\e6.b@9a6(P2EJ,@<TU-a_W:=5g
V:..EAV?.9_WcM,JK6?OY-ccNe@5c8;+DY-7DP+=B2=^+Qe#XVf?2B>4@fa(WOBQ
:IXe8f?JVR^GEDDdB5Jg7dPgI/LWZLL,)?R2G[7d8M&[=VEd>e;=E(Y@DM9(U2X2
LDV+QVOU.P6_Ia,g.a5-@G(>?IG>G)P@/[9Td7/M5ge@A?DU,bW3\>R?Raa=NfNM
.K\eL2BL6:FN9:H6B/W^C.04,-ZQ[CKN:c<3@6c1H_/+=T4c)R7XY87/5#G>,05#
(,EJ6B:QI+5aWS.3LB(^K/R9IXL;O^A?7\ReQ<c@gKU6D^1Q6aYR/GY//(@59QR8
c4<d25ZFNG3(a1GfKG)53cJY.dfb>M7aV@.Kc\_H<1;5T[RU>>-DV8M3MKWNb>\8
XMbaDYTGUDBNO^=^.)NdLIZH9(OS0eTSBNT_5=0<eAIM>+-7HL8M;#4+S&#.K.#&
ZX<M0QG^/GP.bEcQG=29:AGU=F)?B[K9),8:L1gK=;IJND,,QBU=68<]=J[3Z3g>
1=+9;7FTS4/HC+\N[U7P>B&_B>cT<14)#,D/NM\E&7AS;YM-OIVZ-e?.P1WcDS_4
Z:Mb0Z;&\+3S_UERGGD66T,CaH]6DL0&Ig5\5O&L<6/=7XCHDEGP9A0I&&b:>GFJ
W;KTYb+?d7K/a3d#+RR8OH\N#NP7TZ+[OQJ.3LZ(Q(O-1P\MQ_P^<WfA)S1K8fca
3?X?a@H&\CMfbANTJE+433,B[UI@YN6DMMQXBH(VYPCV:>eZ(;1X-AFI7PfbP\bf
C2C-d34B6,3KGaQ^Cc?He#(N.?d??>WC9,GT<V06Y7.^0?6&,a-CLb+M_bQ0@f6F
SP<NEW<eI/+.CTCC=F;\8#Z71Z:;.[KXU3#@K;J&_c7Q.YB)F[J+>ZdGDIO\LSc:
SNI\60\W&IPB>12_B7=R7c&C:]>/)E3ABfdEEe_aW^FQ61GG]c[K:2N,W#^3^V>9
U4D(?CTRU@A_/IE0b<\L45.b13g))(\P.fIKb36M=Z1PJ;cOJFW\9ef=2C<ASB12
dOBeDO986[V+DZK.[2[/a0J+P5(>(E.7WE5<4e(E-H)g.YXN96Y<Y(^2#/KM8f#g
ca#Na#W8?0B/KBU9Y,g>X8a;<:6H2/S._17g-_39BMI)Jc;EWJ.=fMU#9R?RE(//
:(;e1Mf;A7M/AME,Md:?MKST;J&e)-ORR9_(J61B;=W^/ATV95+;d)PGB3N.,JL(
L1PaU1@]dgg:_UdE@dB28YHIJV-:67)1U+>AVTB7#U8.@2&J8MFU.81_\cRQ1+0<
9HNdRL]LTV]87?E+UTNN=\3^=ORO3]_f?_2N\AU>c&?B6_Qa5DD9I5e+XKDcZLaW
]:g\;dT[VY5E?2_6#GWg/&IdR9LWDD_[WdK-1AU/Yc@QZ#gR7JQ?OKO28c[;>f2]
Zc&E>#6Z2YV;O9_NeASZ,W@=1@9fOad=JCdbGSSa=&MCUK.0P#ObI(#fPcLa.d<Z
dSR/J#?[N+LG-HL(EY\NUPd1IM_VD&NeD\C[5T(3Z1NS(1UD,Fbb[fZaeQ2J:dVL
KBY&1I[IOae\d)F-f&e40GXF5\LHMM64d)fO]0MT/VGeTW\f.M01PcP3KWWCeaS:
OWZF-I[e&dJfIIZ2031JMG^XHA;&b(UDGbLNR^.J3Ue0dBZbITX7=e;XJ?A>e75\
F4\g=S;H_cS)._R4,2D^6FF</>UaYcQVIDBZ7NJ,]/X/-\0:IR>8&fM_F@,H/-PO
]^8:gGF=D=2,6.^LU(M0FZVPQZO0Z,P_N)&AGQ0SZDE]B-4IVB6Y6+K4M^?I2Y7P
S1D0HW..5YHg4O+[SF[.[M(>fU0)?)9K01Q(MQK950IYQI1@>bDUU0)ST1KGU_)#
(6NNA^\I&gfbF.&[KT5>J;S:O:U;^E32#-DF/QG6I;.W0a=#K<LT_1\G0Gg^\XS\
=3#JKN]R:RdWFF[GH&TSbg/T69N-(cU5O9=Fa^@DU/P\&W5SIHV]R^>e^X5]3T2d
(e5U<3F8=.V9./P.DJ&>,DaL[f^I.RD\&gg)O7P0#+YHX-Z8PE=G^T.79V\[,LWe
<R[Z]a)_F_A/(J&Y8M^e=+DR,(J-QB\077aKS1XK&DE7\WUGae^5\R4M@=fWGFfK
LBT62VW;&f<bW_Z#9gN+9,Jd(^U3\W5e8,bIL1fg(,<MHcQR\KbT8YGNa@(b)9Z.
19V^#Qe02BPJRc7IA[P\7:V-8&^c1;L;Gf]d(<GeJ<EY>EP#B(6A1Q(;\:^e>^>O
DKI[?(\O+J1bFJdYXP(Z4VdaYPDJJScf);P,Ye?7YaBRT337Fb,cGE47M/@\^T0?
/[g87Y9R[,GZd#JTT@Xfb8+.OAU\&+>0a4:YOAVV3HMS^N8fC\^;b?HOI2=e>?Tg
I(V7(D2D7-b5\FJ0f&RgXbJ9DRD3,I#,c:I7VO,4?S=M2(&g137<_fM=,5&ca\+N
W?:UEVQFa4Sd-_\CK_9b\3CH__]=M&0IfG&>>Ug-@b4BB9-Z8;._?2ZS9KgC_c35
7M#9FOM-^fGF&C<Qe#N/AL0X\>=#;CU]]&@,/^4gNMQeb^8[XO,8bK_U[[-^gBL.
@8_0>V_5+RZ_7a-77<+<I-EYAI9EZ0T/bS(8gXGfDeQR2g4H?=A5((AH5G8Fea;T
EfET99aH2JNDAP;7,6NW\>3C4B.ZTf2@(F=,/TP1cQ0cb3S:7R?X(<>@;AS2/32G
VCS39F18A>IF;<(^eK\@JZ+(QX]9\N?YGLXL5dQc>1@NXSdSeJ6;MB>;O1_@G5>P
-e;TJMJ:[N:]=J9(bg^[>1@7.RNKb-F4KYA]c><F1,#XZ2#He63LG_N=RLS.g@??
IG031J.^X^@?M2Le[UY&I-EPWZ\0Xc6a=KDNP@I;?LaIcA1G8,HOa=)LL#Web:]7
MS.)CgAFa;-GKN02\APMP#IMM2FX2LN9AA43<bO:.;?9OJ;5&F99@?ZQA]JagLIZ
#,+,f8/,H=C_00-(^QcaBF<WQIg.7.8BABBRYS3aUgAPQ@UW<T=58TddUP;J;78T
@-0CLWW@T)dY1gZNROTPf-3ZNG>/O+^OA6_50Ia@KfHL9E(40G7b29<DfM,E:KE?
fgA8OPP6I0Y6W&4S]4Y4-IIOI?(;@U@3E22P1EgS@O.O)_dLBgf_K#d3Q<b7YIIJ
HO[b<Y8-Sd+?NJW=L_;1.1<GYR8KaQ0/cZISSH#C504,KAEcObY7T+]I/H\D,:;D
M4/eg6SGJIe[OQ2RW<0;T-IP<5?AE&P7]3:&bW4_H;S-X7<G48>0MSSB6C5aC()S
X;?J=eX(R&Ea<Zc3M/@BG=<CX7,/=CQ6?0f8WfPG1WMa]N/S/cd2B),ZD)XCFEJg
fEY4=4e\f.,=^>_[:9gf69X?UP4bE@Cd1^TGZNFMa+cH\AM&4C39TP5aR<7R^_6T
cSU/+P[W/>N[Y\#fMI6Ja_H<@I8?Dba;\<Q#9.ZEN+Df09^\=aFCeM(X#JPf<C:d
,bB)Yb;T<,WFQRB4^1P4SZ@S]GW9<XGOecF3W32SSA^]@.3Ec8ORAM48D4(Re\1[
N_F+V?PYF8/8fObA@+E26Y71ff;3f/VGJ9K4<LCcJa3Q.R;f2>IH6:N-_U2e?I.a
<PL2H_eb(.EOb1I05IU02QZ]\3T^#/1g5;]gL1(_McY&OHdR26g;UVJ9HPE]0b82
S<8YD;VG]R9If#4Rf-e27N0gD;W#\A22M\4(Gg[HS[R9.X,A.,KBUBG+3I.4=VWM
(=F?_.9:2#^_:G?JO:YRd?BO9bTCaaN,Z))PF4ZNdOX/\d=VMEV77P4[R>4<Q42N
<a@S>P8&+>K>Z7,6<UV]FN_AXIPISF=;,<cA<dR(U6HIQA#TNcQ5gX.,ge(_M:8<
VO:e0CC9c4R0=6HE>MJ]+<4\><I#VL6NXZ)\MM7&C;4?+G_F6E_<(D>:U6WUAJ5U
gH1M57(\+<[A9:e09B0O2@)EN;^4f)Q.EF=2b9F]^[W?T8.4:)SK.;L:O-1?7CS(
S0:UX1a3b?<N(^\TL,J>3+[g>O2XO>K@BaR81^RRH1=S7#Ke/U3(K.P7>7J5Ng6T
=;DSI@,+I;2efBK9F0656=#6>X?5e^K?3;T/+f4M&,W?.,+^0a<g&6MQc2H_>b:3
YMIP32SZ5DaTG0Oea;@fRQN<T5K:_YL7O888SO2]7\+>f\IDOYZCH,=0QV(XA/CD
,#],&M>f-8J5+129gJ1^K],c.V;.&,H@(/^ggcaCOD1?))gJ,YS]VXO-Wd:1]A8b
&]USJ);ae0ZC7cfY-=?I=(5LQOV>.W1OaYNHae&R;O+0e[,cG&HA3+=X116.AI.F
V:617Z9bOA+,cREN75LGMAM\)]gVWV=KGQ9VKVCR:gg#S[UR,.\>dY-;>2:GY;Ac
KY(TO.c_X5>N8?_2(\JeA6T2e#<E-QFcG[VU]Z)X.-SG8R=YLEK@R7-f.(]QTV]7
/92P;9\]EOJ&>c&N#ddDBAZ;CFJAC5T@NLHfa:B6:JYWV-^LL2]XEPXY+(F_Q9<5
:>7?+XKYP@5[.4_1c2<H?M54@R.Z#I:\=[+<&UEG)D4W1SW1WBZ<W>7B?90X[F5U
+Tf1U)GPHL(1:Q/bI@))<7E7XPZ:L/<SNgZ@X4Je0SSAD<(:G=&-FBX+&@XQF:G1
Z)1Q^NWWPK/A<-H]MA3PB<ER5PQZ\E_U2@&CM_)</)NCW3Y6AL/F#<13APESC8-E
>C@D2)IG7L3)GgASBeGO<-<L<dK+cFZAIb@?\#M^<eW_FW,EAfMKX#<Z8.EUPF<8
cIaG-M(DR,<Y>D#QY)eN4Jb@8HbI,(&ZeUL12>Y6d?&bOdCcI4eabU]?0F4<I?9b
6(16aK.g.P@+F3K2?4M[XUQ@QTN[C+<e?A8DJ-EE+IK]GD5UP20[Fd)fY,V1_E7S
09C4/P>4QHPK3#Nd6M&(0V+3-GNG7e2TB9(0BMH]OCRIEXQb)O7e1RNW-GZ/MICY
5:/<M.Na=K_3-<c/^VL;#K:QI,gSY<ZI1ZR:\27Zf4=YZZ_?+TJPbQ4e2@V95IMW
1#G&>]O/@S5a\=_[[aB8cM[HJGEHbRNL-9e8;?g/(.IERd]NU\W_,78Lf&PIV8CR
A+aWZBX&P.+C(U7H][9XMaIC[B-gP7IQ]S[;NWUNVLgW;O4X:S1@&.]EEBYL58-0
Rc:g648\:J@bNXA@XJ&/C=V,00PO8)H(0X#.MN#IW;^-Ffd[.+SbD[TS,0@:BU1?
P:_?3:<>2P7SM>0K,?:+=.\EN?D9-]IY,F4IHb[)\PD-(3UH]4;IE;f6+_8(FT+5
8#_b1:N-@YLV1ae+IVWXPW8#A(eM^cV&O&#I=\cN5@fgG,S^E8NMbE\b50f3ZF[a
H<JdKfF5[.2)_/g\#[D[7HZ2c&RC67dg<[71b/2CWA_)Bg/+>6:7B=.K_4JF)/L@
3b-L\bN&+E#fE2:F/gUU<^40B=ED#J)HFgObOU3Z)F@\)O_&S8b539XfVMPWK=4J
M[RcZ6.&GAQXbKQ#&M7=)^[4ACCL;UX2664OR7[SRL3dC\/(CI_>XI11L#BOA(4M
DP\&0JbaK5KZeNCX(YDf<(GSVGH0CUJ>Z3X?+=2B.,S\HTZFUa8Wd:+M(EKHY,,?
aT5XHW-;Ob?4fb76Y2JQ.<TG.5/N[3IAWX@9V]^LI95c1TD0,T([N,NSPU^&5RDF
b>)A;CX?g0:@[Q;]G_AW9T3Y#deW=c\.@]Ac7&:?.fEYK:.R=([Ob-H=>V+Z\4(<
8aPd\/V]&2U<PBC)3UPJWJTKQ0QAM=[6ed/[3e&9Y8WKG^G&L9XL;A_DY62C5&X>
Xd-Q0SIK2W((K5SXY@5_]gUOde9&8)PR<)B2<387VV6M_<>P\,GH0ee?O_FP\SY@
Y_g8YfL179FfEE<4+EO:8/44YX@5<R&Pa:35>:+;gb[5Xf\E&X1(]I_Xadf8YIGF
DLgO70S&e([REa<KaOeJ=aR8,<[N0>I_\(LVJ42ZHHR?0_cA@cD>62YPNXHW]g37
AHZc-a#A3M)8NG3FJOQRY>S>2bWINOEO=1+LeQ=TQOc7M^J_Y,K7^N=]bWZ4[E;E
J175EbbM1XYZPf&7)_Y,X)=MGQgcc?cC(ATQWgWGgD_4b->?<[8NdgX=U-c+36[K
@eNLb.,_=J0e<<3,[,<)-Ee;SW0FPEXFFZZ[M-d<UFF06Kg]RA8=dKgP?fXbX<EM
ZBXgQ8E?)(]MQUX^(K#U&4IE]Q-efHOA#H;7T-3<:1.a2NJ<e+OYSRL>Q0]E9?S#
Y6dKQ&SJ&FT:;CMbX0K+W5@R=1M&e>ZR0dD.f@C=X.FOILZ96A;E26b[.@#&g:+R
dKE.AJ-QAEO\)T1Z[27bFH_D#0RAA1AMBKTKT7/aW.AG\I@5\)Y8OE);W3,NXFR3
T9&D3MQH:VLNGP1I6);C07BAc3P:WT6-Y\[(_QVT_+3:+g<CDdR2gF8=Ha50Y)C1
;^6(DLf&G?GX5+BY3XPBUGfOK-[Q>e;>Fb9X7?:7S1YaJHb=2gACG.8g;V&/I=-b
-#UJM0>EQ&\B+N\7SB.6F]b>S)^,bb-dK,3U&923;H)1O/]0(1F<X@CaAJ]15A]8
+OQaO&:#6J6GXJ.gLK71;QTKBOLfQObKH7:cAR?J@2V30Z/<7T/FFISd6T+^3MJ3
F(c&)VW#KfORY-68&cF]0C9\WI5[0.O,g(G[BaVN[JZ@-TOB&K3g9&fGH)GdbBP[
SHFbJC^3GQ:KI0#/L5,Y)K=/QM&=LD,26+C+J>PSd/QJ>aAZ:gFW?4A\01D3+Wa-
L3(=,FCX..:.+J&E=T#GBGZ59C10UC2<;3CZLBbS+O6<RM17D&WGSK]I\)cb7+52
T1BTFXWI:<#X40(\dS5&eO4<O(90>f<:KF4U)BO><BFDZ5-&N#A7fIE4-ON+)MQW
d.^&)[@YGbdd@1_U8Kd5T^0P/7&]1FQ#DNB,9b86L>[5DeI(&O-TDFV8Df?5[D?_
?^KaOI2D)-Z&G_M[WF#S^(+@e#X-64#?1=QV<Y&.eSMA^+K-MA]^C#XZc@NI:NQB
@LU:9aab,]?dR&C&L\B^<6R.M16HZT]dbIAN/;5IV^T<-A+[e7dB8KK.HKgG.RKN
1.>CO;#>3I9EVSg>7b4.-c;/P(=)YE<V,Lba]/P3YSYG@U8@7dRG([SXMR9]1)_C
7,0O[#-2KB41Zf0=E?[?;SE._a@8J#O;PeRQ>@39g4@aH+73GJ#25cV\W3OSHX^M
X/K<53XFf-CT@a;/d?^35>LdBc2gH5_dH#5I5>AU/37[-C4EG8;<)XW/9OTVD^/)
]>/VYFbF_>TG+f.3WUG#5=QY4W37@IQ5B.S,5KH7CG[e.UeVCF/#S?]N@]#P>bE5
<I?C1/0HTM+_fGAFOJ(XHfHER,/DOR>F9S8O/4E=2PTDE80]:a:&Z,H=Q0?P.BVJ
IfXV):I5dEI),(?5UJ#be/\>4;3/\#.&AaI6,KM0[31V/EUXEcLee^/JV00X8NMQ
Mg#K\Q)HGd<]9c[77L&G=1#K-?cWb.9.e:JTd0T.IKJaXVDALaPSCHO7-J\Ze]JE
WF_R9a2?9W),a@DKB5S-75(TK0AgZ\FIBSV>9J7>?XOL7_^JF)1Q4MW9-#;X<DF/
2U(Oc,AY+T?b.])>/[WacJ;VTKNLO:5cNI50IIJ3+/83E=?@cc:LS\Ja0(505OUK
OB,H>?a57dZ=IGJ4Z:B&W;,EXXGSBIf[d,B6)HLU<aMVFN.&?SDN6K9J2V]/X:ST
)WY[>>Ae])SB6^1JfUFb^:HC1d3\bf/]^BD&UNXHTb=V0/;ZBS.Gf^aNPLF:3fN&
:K=N0CE)/-60]M&B-E3;\VQ&+H?V[:(7a)c,JH5>9,)+H&S<&=d)BG&fA6<_@E7G
QfCJ<675/e>JDE8E67>WDcWTGac=U\LaUDNN9f+U@R=bQGJ@La,H3P9g85,Qd2>b
OgZFP?a]5PUCUVIKe;=7[H6cB>IW_cI9FXaONT<UA<aT\T#IO.KRe&A-N7R_IB86
&eQT-9M-6(]<KUaX2/TG(UR&S?&[_:S]=;3<3+J&#9<)&M/FgC@:c75Y9ZYDQ2D4
,OL;af/R6.,[-U4ZZ8cY/?;cAg^8JOA[Z:Sg@]G([:6TC#HGVZJBL\\DLe4)+T:\
Hg.@W[XNaa;:bFcBTWMQ=Z=^ZE:;J]L+1_I3e6R@2Q./,<_:JU_-Q7L[UbCE_\-b
d5];C9c&c5g,:66_0-0CF8_A/AX-@KWIaJW,E+9dO5P=J>\9Ef0g7OVG,^,V6.]@
F8T9](E5D#QaAR:<.bA/6OXM=.<aHC@5)?-L0V?2M+g]R5eRHNc@Y3RYZ4P1KP2.
2]/5),WL0,>SBf[1)OIW0.Mb(8-PG@[M>f5BO7e0a3)FB)Qa@TXNV6X2G68aF0O+
9R4H[=AA4;cZLF>/([IBA,,(IX#W&8dCEE[R?c-9Z<1F+09Z0Y9;\K<SHT5UW.EV
@W3<A/+d#4MM[ELbZ9N(0)ISgQJf)N0P6^E10^4#8K4YQWe@d(.bbD#S-<TMJW)_
-XLf@;YbWQ#C8CAB4Ze4.?>3QRH3eTT+XfO4Z=;,SF[PVKQ?\PT8Z7g?HMZN@)^O
F)72[2)eE6eWM@f];G5[gS(7F3>ODR,NZL3I\>c9@6&KL+F4GSea,LHa:7?+G2Pd
IN,&D>,B=#_/0F8@M66)ES5H;J-]+SF+/ReAL\b4LO@eS.NN15;bga5R82Ia(0.C
YbYMTedTYO[4NaBI^;;d=]4=,&fKS)YQM9^1P-RG0Y&Va1e^d>53M=@V4>R89KVL
dN_D@=@<<W9&M6UJ_R.36Eg?E#?I9]AKHS4<?<8f^)MQ(,:ggaX#V_@9TE\YO+R&
<Ua),[=[]B0[1NDR8USc^&L5.?Of3bWZdMf6#\BId_--^.5Q5fK6OT,UZ/SXIY16
WL8<S:]NE,G^2XG6K4ME+.B;PO6ZR5[[8V_d7QG/#fMXBV;6(cSR?dGb><N@a<1d
:K0g?E:Scf,2aM2KXTTK+GCFCBO4G+<LN2DE5M[?62(B;MFJ0VD2\3;(\XBRIW^,
Q^V4XYA40Dff26V@eL@cYE6/^XcQB],13BXTS7]:KcYb=2WL3[,BB?6OX2BS;986
)e2=,V854Og]a3Y@AN(6HEB<8FOW@a8,X0dEg4X@07BHKFC60b86G39>32fD:HB]
J_C#7F_+2MCV]NL6-8cS]\,M7<dBZK^8Z+5c3dD&_<<#V:&Y#dMK,2ISS+FK?_1g
[1\e38EZ;NHH]?7-K0aFW2d#fW)KVb_(5-9/H;M0TMM70[7:D)C2RSHb7ZF/<)T0
Jc[]dS:SN_MFP+<L^7d7Z(T;.2G6C([7<Q<;1>cXTR;,L_bTgO3AcL-?6cN6KI[T
@84_;JA>[KM#9bM8fZ5g]@^0UQBT>QDVTcIA7J02bTcL_O#<D>.+;XO+(6KP?\Hf
@7YR]g(/WWC9)+Y&_/=FT#^JB&9<b[E<P@JX#e4&PF2<+KIV?=I^+S_SB7V(Q2<C
Ne(#0.(U.d7(Y_\H,SQ=OZ#a[;G&_b+=+30+(;HTOV?/JN6Y75FO;.<G\3f,M+=g
JD\N,H]fTC3Pf]=;GD)EQ/H<@_YcY@)Qfag;R_a7\?D^#0(F_d?TJOK]5=<C2e>Z
dAc/:ZM>Q]U<)6WeRS\E3.J29a-F4S6V31SI^B0U73gY9_=LJ^\.M#>b5:Y5GPBD
PbZDD30-C31f92gWCMPZUB]XT/Z]SLc#1M8T8C-IL@M+/e?b\O8RbZN5?eYF2KaV
VI/RWL>7+d]XeR_:G3Dg-VM.X;>1,9SLW&\W+dG_KM>,?TUdPL7V<aL#LR]_=R3K
V3=]cX2>P-Oa]+H)?DT82/gc)&f<S#G4725Rf]U-/WJCfeTFCQf>O0cVbES]3?00
H:BJ1@QSMHeCYXcIDOb46J9/WV8E29ZW18gg3ST.,:QeKAUJ8>dAM_D,Q:4EXO/0
?FU5X0c9aJdA9VG4Q6/DH\d4+@eX\@f/K@NeOASgEb<5EZ?RaQ<IO4KIf<Q+J[/[
EcCQ_GdCC09f<5HWLUdB<F[+:B^K0;>;P(ZX7a,;WKGC>5);NAZ#>:)GbTV9;RG5
4G?45-,FQ9c[&/L8A[O?3G-8>1e;eJ==d[96?1^P7BF4;6G5Wg;-\W3dD\CR<.f.
QL-+J-X7890?/dUOfG,3D4<?^0YU?UZfdT9]##d>,NB5BA;-eFGNP>]f>MPGC7.T
M,Ya=(KK6YN,&VR9X5Qd+85X(9SH0g)GB0Ug0MO&;ADgb.&Xf>@e+>e@6BFTIL@a
ZCU83?-/CA?@^<[NY\gXM?_@gHWGbLVU>Tc@=GcgP^>2(AW;I\VCFRZS2W469P;Q
<@TEE:,?3=D_g:/E/#,J.D^+S_+CJ12<QfVXDd4cIa6M@OGFSRfU_K577Ia/O;[^
fa]]<I^/6+75gCD6eU&^BSRS+K;(ZTaT.(S;VQ#,EOe417=;:H5VFS&X#X/A(WXc
S/7]O?AUg6XN=3-@6VefRP\^2&@KS,S_<-DL]_^a:RJO49cYEHAPO1?7E-I=AfX<
VJ]NEQGL_:J\SVU.fe:C8AddKVLQ,VR^_eRESP][+6&d\7(M3Tc218]6a(IE=+(H
aQaU:F3I?+a+LL9EfNb<B=B3cY-(XS+J&X]^B5.^:&K(ESPB8N8\R&PAJHDegMG#
5[1#/[1CU_b)=1C#:Hc;LU7@S9M6_a5/B7:1\e)e,UWD+S)[<AM(ag<M=eMg&2aD
G073-3#</07-O<@&1bUYcT;(PZEg7N+^JO-JJA#B3:g_Yg>XZP[9Pc_MI>7:^Gb-
RI^e)OB<JagUfHNaA(b-?:_-QOR6@/G?@^CI);;PQJ\N=X9bBP@Se)4F[YALC26c
-EX]S\L=H.&2D.3=WDH65KCf6Pa1RE#>#X@#MgAc&T.4W>0D-,[[)_;,gaEOeY;@
SSNEQbMQaX<XT2N41UYP40a-.7([eWH2>ZT8QX7;BGgP8>P)1P_1OZccd:C7(9Tb
36/,2;ObWWEUO\N+YEB;.YAVB=_1DS=OV6-^@#Nc151Kb1PV.8?)E78</_=)0&dK
#),Z/W&MgNI=>YI3OdVd>^\@D0X7/WY_JEC1/]SXBTdB]8&^4ZP:<^]PeP0-eR5J
[g1R\d,da4.fCYQN8MR[4gS(<fL1dH4a<0Y7beG.^EACA,T@V\-9KPK:8Y?E24#R
?:P#&GEfQZ.9WT3b#YfVW=c@^,SW_FGb;cQC-,QD9a9Pb5Q(G.fWg-3,1[<A<)aD
e\JA#3F3bQeR^,W;P-bS+U5PVT)92W9cG35LI;KAOKKV6@21_.0+f@Q]f?Z+F=Pg
U;6B[[5(X:F8/5Gg&4)#W?YM]bN?[MQ2bLJ-C0RS.;-Ga[17DS0=O)L<;fB_W/6-
a.?M5[Z@H.C19D2:a4XS+1TKM<4.#B.[QcUG8M=B:#A[8d#CU=TLbIfAYYZ0QH9F
=EZ;&Q(GY(P[ePO8+aS.7[(T7=N:.D:M<>0(V</M0UYKc<Q30H12ZAe?:/JJ=IeC
Yd]JcfM@(C7U6@L;Ub2(QZ36,(O59KQ&B@&:;^PYfA+-S[4+B_Y,7?&X.&ZJ(a2-
#.]3S[GeJ,Z0Fg10;;MICa^H+;]98V\XP@MAB(P_-[Yca?A.?.3)_gCV<C2[W-<.
>?H3>[8L.gIa^?#TYfGH<L99TGUB-HEZ5FW2Ue():f3;bKY:b:):_C0QDO,\<QHB
[0]Z98+;I2[\/U-]IbCg/&eHgN+<Q-;e;aPHS\@U4UJ-Y(4XUNceV7O^]_35Z#W&
.cE#6,O1X7W@\e?R/D6:#=#>F@/=&-Fa];62/<CS7S>d]:XVdN(C<ZK\8MGAA2Y#
@CJ4gJdHGO1-egB3DZA3,&VFS2Y:##0IeZN-_7#c2e=#,5gK<=P01DXS/TKUXF[2
M:HRK=MeRLDA7b(#T30,MT?5fNJ=:RI=<EFZFacAW94+V@d1SYegKNF#G#/T16G)
=2f6^[<B4:(M]98KZL8X+S:XR:)6M&JIX/\OP393EQ.H7E5F7A^g[8#Z(\&(7UaA
+f_Q^JN9SA29ACX;<4#c@dR.AC_0#CG4?8g#5O0eaM=V5(&,?YJDX?@C,G+DQ&;W
LLKg-^W[6U=YJL96,0<^/P-YJ=FM\?2MbcGg;]T8-^>]53L@OHJM+F#MPJ;5YE;[
&gX1dFM=15RaJg6VbJF##\W?GV7+PU7DD.])+)60<_a-_&+5G23SKM0I28Kc_F1V
.ZJCZM.^-ZCV1)9)(gG@3XX@=c^ZZc^\:6\]X;ILGP6<0Z1)H^Pc_WE<7.JUB/K\
8;XRgD((4T_b9G3]]YX+T3CJgI1YSK^@fc?J[@L<ef51;>]QJ_Q6VD.S;8R@DW>L
5@)JR;FUZR5:&K)&CTZXDON,6SPg&=Q=X-FB>d_]gK,.aXXLd-Ig<PGK7/-:=H=S
J8K(-E+/Pb=#.)4+=[FXC]C]6V8[]OJ@=4b@dD^2MWM8&fKW(S@C8)2V0T_-Y/?X
/beE7)f<E;90QNFY;RMRZ5P-_WVWYfIe0D;F91^Q:#S4I3/gZR)YaEM&RXZ&c4aX
Z[^J:=;SMe]RQPDZ28HVO3@,CfFRf[9K<ANF9+IaEBO.O\TN;(#JbJe-5_?G)5,X
2IFRSWLJ?MJ(I;A1,bC+V-M;S(g_6C?AU9,fY-:49/M1_:UU=,bCPcWQ#66---1^
U>@[^TUE5-VEA;TKGf[caPXRK(ANF+&@MO#86HJ2MV7@b?dLP1^DV8+./&B8GPH&
:3gFb\\W^:-Y1<b&^<-Y+)#b8K7N+B\,c\gP>M\S\D(EJM?KD/AL3/)&b?F.>-CQ
\]f7:PSY,<H>34.N&Z8LMNK<T-bgS>TcS@4KK>YO</ZE\Z(K:V48Na=FA5_1)0Te
geK_5JC2gK\B?XL@e:WMB6U80R/.V88=+?2/+4/A)JPbQQDO.K/KQ)A6=.dbAa;9
<R5/c,=Xd\HAHD7XdA,:,Wb_b>V#R2Rc#MRa)AYD4=V?-)]-T]7eL(/-\3aXKSI#
<.H5HD;D)W&J2_I6DI#Z/#+\YPU+6e7dJ,\f>^?4FeHX+?F+R?FNPbf?34ZN/W[]
]BW0W7(Q]K@HPaT,)_D@6_[9CN-,UNN,=Jd83@ND);DF.Df:P6WKN/NMVLY9N_;[
?TW5[.RN#^I6_N6(;F+,HCfB\X+;f8b(_Y]M0T\b?b0@g/UF]GgOf=cF&]#==H4/
F[YF0/Q3&ac3Y9/9f-/VDSBT4@UMP-3BZ/7]g]f?fF5ZcK+9.78N4/(b<JJKb6G,
P@B==(?R_/8KeZTUU\5W+f7FAe@4BE(;U/,#EI\[Of+Z_8EF117SAc#^P2Of1f=4
3691[7([;IgR1P?[@IHg)?_D&2JU6^L.+3PK/TY@WYX2.f9bR@0+X9=fOV=@;eH.
KD#EUM^BU)=fH:AaB6FUOA&IXWJa[U[9f)35S<g72a7Q,^/NNC\<,fGfG:JWGP6S
f)#L^e3=(LE[acTOI-bTN1/;8aE[022c+&-C.>3YJ8>HRVGIK]e/6II^X7K^MZJ7
S0=a13:(SD4G0K@,:HeJ^7T4&0G6Q>9:5TDa]+6;-.@L>3>KbMc(:_YG50F;ZJ3d
/Nf_8BH6JgN_BTF<:FMWZM4<d&69-93O+QdIK=]+C6E/ITWGN(OK/M+e#?X8NN@=
^(_3M4)B2eV;cZ#ScfKeG,8SX9eYED2N..dG-1WW^Y\@?=JW7V>86E1C5(-Fd[f6
031F?1/C]UD#8R?&8H7(eAVd03KQ?/e+YX#OY;fSNg8c2?WDe(&BQTU9G1=<d#9F
06e1W1<F?^A_d7dG@6^BG;+OYO0fQacgMW1DCF1&,:dUE,:b/NeDXQG)AKBMD2/3
V&_5>\VH]2BdVJ<bEW5:5+f5G(:GYV+BL<.YPY^MCf#CIRa2ZYeaVbO)V^^B0>N_
UBCg,&?O8KZ)U>ae1Y_=E+9R5R<a@JMcOWe<[087d2c?V26\;?C>N)B#TLU8=9f+
4I+SN-V[-K@@M,+)]EcOW1H?N<2S4_9<FX06Kd,8bCNU-K^=ccN_fRA?Og]c-Gdd
+G\=DP/I(DL4(O[>gFgU@E2GW7]\_c@gOZ4,7OC:/;ITPMZH-.<)b6ZKM75T<KJ?
]T;<dTC4AgJ)aff&-;/-CaWC(:PUV(3b2Q^S4[M=4.gfIe95HS.>dZfa8g(]7)KC
)-6L?]dLV,a@P;I25f96D2fKFBIB_[@A&_-]HeU=<(&[RPD4C.6UWXNRd7EST&SF
&Z[4<B-XDDGFF&f@-0,8GZ>e2(aJXW8D?-NKFYP;B=57_?ESPT+fL?98VOG75PEa
8f[(O#KHNaZ./_cA<EC#EJFPNb_@fV/@_EPGTV\f#;bVJZ_0N83?_N6,3ZY:ga)<
16NFV=P1OYJaP3^(J&63P<]Y6\GH7.K47HfgV1>,\@SVT.M;\+d9DE1P9&Q(1_._
,8I-L2^K^<,;HETgX7UW.J\DS\Q;S[d/c.cfe#LPT7fN3DN@B>MU/BST,Q__>g\9
>Q-&A#dH5@>;F>DH[4^PSa\XcJUgHabMgZ](56-=a&2MB;?21=<^94YQNQ>_>1Kg
61ALPeB]5][aY&RcdDL^^CV_TK&ZZ@.eb\DGYSJ(86OP8KWF3]4ARK@4\3#KQ0e;
Zb9(\_[)@8XB?64J#4fV69@\[>9DH278X_VK_-(+cgdMJ5[;G-L,G@VX#\fF[cRI
W6/[?eNf+YS4[I,ZNDO+98AQL77>B[:5S-^?85;S+b15d#[AG]QRRTaX;FY/2&KS
e)0TAV(MR66CEg]eKE[((,^b1/O95.H>VbdRB\[0^M\gE,E>0F81D;4bK_A\X>RU
SHTN&KPNYV.eb-H8ZVd/:CQMW#&R/TfZ8;C2&/?S28aR)QUMGaLCX;JTKc+K-&DI
208<-bcE?)SW#@N]c-1N4_\Ae8;O-4Sa\?D8&XYFR:)T0K_TZ&T5SC1,J)I+J/^Z
e^Q-Va#_?V>1]S/14_(=T5:N&2&6@8>C[@+JT0F<6YDB,46NF;3I8Q=\[B^F1\[W
S?X9D]P9VJ.9C=4O]M;_@5fF#e;XE(,=WNb_VWB=/?Z8ID:VJ.<TVa?;OYa5(Y6X
ERF390J63&dGG3?Ec=L6)I,5^e2c4ZA>Z6QP:P+0G]8Lf=C-O:=:\>NGab:If5(X
?fK3@^^L>AJ>b4gE>eY9(7G,BVIME-SI]]P0Q+[Y?IdB3P/,X..OR_D?#&3=De:0
]WWW]T1_5]936&WRa3)fC@cDO5dQXSaXA+/3e#/DKLZQ7UEb6P\Z#]NA]AYJ?gfM
fX;Vb,Ug43Q<9<=G2f2N,@G(S_3?5gSD[[_VLB[),Ve09O(.8/c1&/4A=TWQE#9G
WgU/Zd?:^)fIE8])32\d_b<?=LI[=^J3>94@@EIf5+>3O;(G[V_8C6;4cL)d0ZI>
6c2QXe9Ae<Qf=;1^^NbS+1QcIO6++:AT(Fgf;=0UV3^I3M/f&MOR^PNV<C;G5Y5<
D+(0S.<60Q^cYEN\RX&ZPO+C_)1=02JP(Z]\]PUH7<?L;;?,-c[\98/Fe?6<PbY3
I6IWJ,,ERaQGNe-<@H[f8.-K&5ILH/C)J]O;=WP.P(A1<O(@^#L[Za+(5)Sc,,Q<
)Gfb@HST_,gYIYBV&_X<88C_GEOU#()0#W.S;<I<cA9E#;.L,[,T:E\N-NE92:H1
[T;;KTE;[>0=P3R][UCMAP3EFb>/<_<bOf#GSITfOPS2.XHV[b\bBE<2)4fg&P=^
ZN+P:)=aQ_Z/7.Lb/0BPF?[]D=TE5F#&2(/#8@&7+F5C9g)cX[--c2^3((7Y_7+d
CC0D-ORFJ)>#PP/2<HD(]NKS0W(V,^fVI,MB2R6R:4:Y.L8V,MHY/3Rg9K-Ed1T1
YOA\d0GW6:#CR493)VD]HfPP6.RB)49KT.XSXH+P]_I.c):2eZ4Yd>ZSNRV=RJ5,
@AZ[2=)^<.8bTV=\cJA@=d5[30NMU@9@Te0Z0;3[KC7(g;daaTa9BE:OgRT7J1FJ
OOdaE)b<0.0\;P(.@9?-a1Q<;K#BL3]L^dbcc)Vd&5V(5QPLbHVTFbb.ZL)MU>J#
de#VV7bb,PNabc-ca\e(_+/BdM^RDcVFe#:_7]+(01>L:L8eM3&_b9C[Re0b\/F3
Pg[WJ8FM@NJ2;70/X?G\a#/67f/6GV7G7_>@50ZBB;M<P30;.b46aJFOP8(+L<IN
C^D5JS;[&T4T=,K&FCg\A;SSME;8W:M/9M.:9c&dC-PAY)#5?YQ?SL)K\/F]0=WD
.C^X>eR7XRZ3CXVg:=JbU+.-eee02-BgJ6E-D1gBZ(-F.R:TT?):AK,f,+[X,Q6J
J?KI&b>+-3&7dH>-gPERb8.c2.]UHSb5:fO6dYZ]YWI?8]Z+>1&aE06e8-C\FGfG
)5734/U>T&;a0U=&aD[PCZ^UbF:]W>1)fL0G@8.)Z?UYJb2:HU^>FP-CU.IDL^YO
I,g[B[.>:15C2H7;GRW7gU1eM_d1^=HAJ4R)#:.+8]1KA,.?<VZR>b+YP,2Y>13T
XeC]F,Y0<#@&PHD<?1F#D3.afIaGV#5?MbEMQZHI@1&I=]@8eMac(ZdeQEMPOc@e
d76#3F(a[2Z@+:5MUU7)?]_]4+/A<ZUMFM0gC4L,NL=+<J_OJ-NTZ_ZEXOE[Rab@
)#ZWHX6d_3FJ/DG2L5^5KH1P0OR]YXJ^UQW1J1@E)_#LGXDWg:P]]A]14WQGH#T^
9JV3bg5QN8_,N0[57J3DPPZdgA1SG2T/W=29_<L>/J[Q=#\6MC^?aWNH3L[@L?YL
\RGTa4KHT-<85D1@<X+&V0C>[O_b1Vb3S^X48O;HWU[Y>CW?0CC,@JUV<cP6.TFG
^L=A_K&g+F8S^f)BC@K-Of+D:DNY>P=I?a[/=[<g:@T>JW/T\A/,CU^_HBIOf)E?
CR)+Y+B+;:],E4R<U^_+fA8;#E_Z_P_7IQ8.fCQRIRC#4fANYOT,AYb8E-UJ;2ZQ
;U3,aPAe;EM-\DY13U:d7LLgNIM#RWF\K\V+R\&Xe5?_8A6a.C9M9X,,HdI;^<O>
516MFR=faYY9BLLV2CX)#:=51=[>@+C3g-6dE3CTRa13XCIgS:G+10T?V&SUD_H(
A:EV^1:RXVdN+>FUYIbO8B/L6gRU_L#(eJ/J8NQ?O[BZKA<]d8Sf0<OCX.17[Ec&
CG>RPdW\N)_-B<BQB?V]dT\S00Ea4bG5^P?c9_I4[,<,QM1A8/D-8f>M<+Ib#gQ?
:VZE9P,)C&X#J#g[:@V6QQO0GgR&[:ID@GD>)4>7f/8B^46H/#STb9UD+;_18?1V
_0ZR:I@JN>U_XQ2J<Q<]6\eG[&cHLe#V63[:EJbdG@L0V2MQUc.ZJU^OC/XAaV,T
N4>7Jf-\a8F,5?RO&6;E>XSXN1WNTOTc4f,LBF_SZ3FOd<6+K=9#H.LUR@bN&b0/
bETQ[DI2[b0L#:)ELR)8#94H:>U1E#H@[Z\XdJ;AMD\H+A/F3X_V.^Ta^#<5BBFG
gBEcXTg4?\K+ROKfNZKMMg&EO\NJI[0TZ(F0d1>AAZ.a]M4G<LHB6,[;(N@dOO@\
YNgcBI;7A7E@K)6KB=KWaP;GSg[e?TA25[+a#XXCW<]+;5C+NVEUW?:3d.O<\?_S
8gDUZ7B=AScYE02B1,Lfgb@f@7#KUU5bfNT,<HKI6cG.XaDF5E3_bB,-TFFM4E(7
/4DW\cX-N\EeJB?KbX2_Y8[3D.@eV;c-c.)OG:[OIMBb_-/47SUA2DZ83@2TVV4.
O_YbH/V^cFE0g^,YTXUXFe1[-daT@a;/0eQ/U.7NE+5Z8#L<f@cPG:4VJTR]/dfS
((1@dRMN&74E=<6[ZG25Z&-J@.BcE^5Z2=^OMgU6KAG&bOeGb<CbWRe#K+J0f5Q#
2LJP\&Y&<OO=YB76dE>a&5d<AQ[)0GH-EX;DW96?8\0]:^O^VWYe-6+SENT;;Q-J
Q?c^LH&Da8<86BKVEaK789I#4_RA<J_3TZ()JTb[Xa-b7^B0NB[=WNO+CbH(S36?
_N<^@<e3=]@W=FEG+RE<L=O+G_D@)>SKF6S[:.fcA3:#4PE+]^]VS^@P]WFe)cgK
OF1-?Q8)b.P:&V)-BZ1(PTI8d(#1@=))8fF&_E/KXHaQG=^JY^?B8/<MZB5UP@K0
8K0OgdC2.Q;HAF+g0T&g:&G?@e;US8<IP@0W864MAUdN?XN9NM&4@-94>>4@WFE/
&8VUKg5BT60R)KZ4(RA3TJ&3E/H]Q>E;GY/;>.4)C9F5>#KF]+:9<e9c0aO8PQ.1
;I@M1ca-RD:R^eLZ/g_O0]F=^E:[^0gNaJIRAQATH.Y>>J9?B1eV^;15^C@ddN6J
dcN24WA+T?:SN>e@G;B,#3^e&G2DZ=c0<]bC0^dSdXdV\I9TE5Y[<BSOa+G+5.c7
:2&Nc/@cTLND@-c<gYSaG=>\@f9b+VS;6?L50=DBYZMH,L.YW6)?7^S:UUO=U86c
=a3b^V^gI);#RW(992LUCPgY8_DN-#.VPHC@RTA:><1+#&-H?P^I9c7-2FEPfd1O
Z[+QD83PWX;\Ag^-c)_#1_44/ELYJ,5L+AO1YO#,^[SLU#-(]8&73X_G9/DL@9M;
G4Zf9HN&UA]JC^SIUe9-5KPOQ.Qa22)3>/C)/#H[],Ff^[.[KZV/Q8&>99<TSRZ@
:\Re:EM:V:\K@SRDcV#^I&BWE86(;SO5@1TVGTd8)6#_4Qa#/5+[Y<INVZ=ePE(O
=.0ZC;PV1#DV5;DAN\&NNGC+WcBL6E]N.Rd#.84f]cE<XV8&dR@:P,QZ+^eIPT&C
eL-=Q\H#aOAD_&Y:<S4ZaLHLAc[V7b/_,Y(Bf]\;=^:7fC0f5d:&<J<0)]+K3&EP
/)9&CGN)1WBW])#2BQC_8TMfBRSW,U26T./8eTf.=CR&\5[?1ZE+.O#)KbF=DZ<\
(UaS3TS@:a9#WULA>-M@9^Q4Ke6S<,G<S-ebVV(@e9&\c1WeQ\;I<6fTfPNeJF=H
N5HB[G6/N1M-SJfBeE9J33:?0?87A3E=UP+bbMG1OcW3cc2WHWOUS54a-1c;TYK,
,)4[U-?_dHQ;<1(B?g=b[8+f7?IJ(=<57X7XASCQ:?8Z:IVA_Ud.DAT,?UAc@Z2K
dZK9]QbYS>\OJ;_=[)FN21;0P1dFb;&bQgHS,D-K.3Y12?)GZ]H&[^:5,OKL;WX>
R99eZ](_TDd1L[edE<_=@24-5@H#4^;B=cI1/1#(8;HcHL3_,3c\C_a4B>IAdGBT
e9]JM([;@V@BRR_RTg17B/1PCabO-T>OI-K#MO&2)S[d/d&]AU@d)_g?#R/(NQdD
6E8H[Vb1aV6Ra4GIQ;@2R=17g1@-0eWFK-4PE(c#DU]()O[VWX>.KCKeKV4E<?HW
B@:&a3T1Ge,cRW]c]d/(+ge\;J)^BRL6AH-,2eXdGZK9&A1.)]PfBCF&>^=&,Q>/
^G13AgZS9@FfY1_]O<]KV,f72GE67;YaVRGBJGI1#_/S3ab;bg\C?#gI9@aC\+K+
bSV9f^6@]geV^EY.HeXa1=+f-E+4&b^4G6_8f66LO=T:IFS3]FI7XYQZEa91_)+X
H/d\X-XO.g2FQIg^\Z-AEL]94e8CGKKY-B/bTF/#KC+>LEOZC(&;N\XIIdLS#c#c
dOKG^1NVT;eRaWT@.?g]+5\U\:F[f]<>)HK)CE3,LW6[:&&=:EWBW=bADa5?a,G-
_(0U3><fZH3@A:<ZKX,UQE.-FDW_gNK=4C<2Z6EPMN&I?1PJ^S)Y?Y&#WT?I->?_
/ZILJXHe#a<[+<04UA-MfF1e.A;G61c2ZYWZ45JQA7_6#9Gc.#+eG\MOF+5/>]=<
?=#?[dDQ#g;;<UDbX:>=/K:\]+ZXPcK>X=D49-)_5QC+7G<XR^.BA9(6&SH6,1O+
KN9\B=Dg>YReYHHa0^fKG\D+G4-W2c].d[JQVM,:B7B=60@1,gN+(IYS96:2/U_F
9cVAc1N39>CaY0&_8Ne@BMI8SdLBb^>#O,0YE/Q::?QS>ZRA7?+C=&Y@@6YK0VE5
FD0Q(V,IK,U7cE5U>2<ET:_4/(AI/.EHbKTX&N#^SM8@VYRGQg>NVHI2:3YCO,L8
GRH_Q-_N=?Na^L6<S/,2/?2bBI-DKfcVFM[;TdUR5c/]]54Lb7S1G^<<G]SI:FW)
KL;>.Jf<W(P-5RXf9WAHe5]R;\RT;<>MPX+QgS\\f6KE/.78>4d;)7^ee0M8b_0A
]__^R]^B>:9ZN5^]ZJBE#[M#1;@Y039/N>25JK&X)[S,b=6;d8Me[,3J;9BNTTKA
;IN3)8J2I[G22EP^Z.7aTVG9IadGP7Q627.U,A>X7,UT4-9#UF?QJ>-D;8)W=D?d
g<SES88]X;&D(XDY#];>2bQZBHF4BNf6[+)V.)(D@>LW@NTAY88LJOW_g>X)D=>J
=<<B5f=6ASdV;=b6KH3de]=V/L^]XO[gO.Y3e6&[7@aPdc:aca-QFFUb7@83[ZW.
XKfB0&4VS\?ceeC=]]+M1Icc6D\D.#==+,/)V(214F4/)97(NPK1U0Q,VQb)R.DI
a#:>ZAc_5L,W@CX(2W,U@X5U?N9N(,Q]I4GbB[e=NDXUMfQ+0M,O.A;-I:f,LfF+
=2P_)CfLF:A+-,M20]e6/HQ\MVFIGI<>NQ@1@@TMKQY8CXLbHc_SB\&7F\a)?.[4
UN9?5?.f,)YI311]JD;RLAFPdI;&+.A7Ab2^Z.7B?YKZM@)>9/>&;G)?&G\c)NY=
S^TL<F3_-</4B=BXOXG<)CR_I,PbD&Wf4ZB-ZO/DIN?9.aOf2T>eC@cWe__K.U+A
J.RK7-&+82ME].\Y=+g[Xa.gg/77F@^:,#;P+)9-M?//?LNB8c.5L^N9Lgf04:Jf
XSVdD\NKT[G@F+c14\OSQP^BP<M60ME.QE=YDW4:JI].Ra29)\A.]_/Z]83OQ;?=
DV7/S8c2?]+OS7Z/IZ6\V0eBHXQ5>CeR.8dCZ2IXG&;_2,PaHH.;6-N<1Q)F<;15
U?NG04D_6P_LMCa]W-\;>R(.@0AZ.^YKXbP&/-B?P.]O3BVeSJ#(aB/OFS+UQ6L9
TM#M7gY/P#H-3U_YVS.E^Y-HHC^4-+OZ<49fX8]5c3LA\<a6gUHf^bADJ&0YA3<K
KZc_f.@.f4?eX6c)V(NBbCEA:MbM;-T.:BB5=PC0M/=AWRbJ]BgXS;;@];4O.eIf
7JN<_WS4ZcD=#L>[Qa?:-QK(MU(+T\JHE#8eK+^>G2&Td-S[T@BRK^<2_Q](6=_D
F9\LM/C;D:^1bcDfI9^GX2UIY(?HAG^<(6/C)12-PE+N(+H.C9@=G?-B;L/8):c,
N2H3,DA,YWC0?;,+H>C=e#fDIefI..F].^HHLX+5PCN,E\3:<A]:[(1R+)ST2L,7
(<3^DV7+Y(X@BI.W(LX,GJMOUJ>>ON@7>PB91.>UYVRP+D_\95Oc&2:D;]eM]=8A
4).ZNR.THL+X+<J<1BU_WaV,+M77E[@7]KTI7F^E_FJZJ?cT^</CJQX_0L(e&]f1
ZgY_eVGTN<71RZ-4476;CJ#IKf.^6#8gHB=2V9;C/:;[T/eEIWAe?g_A+=M8_E:9
d0+IbAHRc#7&gP8R,7c01\[6&3(5(HD2Nf2AFg)Ad:5>CfMJ-\gC88F2<5<bQ2[P
FY]e2A47EL>Le(XTf5(S\(KQ:S?5B#X^9210<T9RQHI&]B;W^653\)UXO\,CN6=g
GI>eBZCXJ^d_CL&U0JA[NR\H&[UFEBReJ57:PMA,e(5\(+R+Y,YPDXOR^D7R-2<O
DD.RDYI47><KLgXE7RA1[=S<OCcIa#21^\[HK@)IA]8e/T)B3U8f2MQ22U>1];X\
:(S)JOMGIM/B)c]CJ;B@#I9Cb7dg/f6)RLcFeMM4O^]8D>IVXB,=bb5#.#(7>[K_
KeEOa,&0V7-Y91G^5@cLR3eE;3/JE(<5X4BO_??1:?;<>>=72]6d0=^+AZ7CdXe^
X\>3Ffc[\X<(U>f^V&5cS^-&N.]f/(=P,(YKF@_ZbMf?G[4T.IMLGg[M.Y6B;V21
YV6FB;d,:-VHE+0M[cRM[N,M:C<[0GV>MP?CCc4-9BPQbWYH-e>ZM_GUdM@TF8a;
9BbFU,VP-g]fF>RSG+?2,HVe[1/JGN>(IP@87CRWU(.E>N+]:S3229dG#\M80]AY
&?.;#F.D4&cSd:MWAD([BNQ&DV?QCDD6L<ec:0L-Q;W&@ZV^.(X@W7,RC4<a0V70
QPS2G,K\PTg2b#NF_bH4LJ)K]W4P(UO1Z2-W^GTO\LeHMHa;.YX2X[dc-S@CZGId
;IRU9g>@_F-J17+.,eD>-]_RaI;W^c@&COX:EH?+NSeccFM;d3RX.@AMZc>LIX,@
OfXAD7[c1T?E:R-E<Q6VZD@ULZ6P<72V1_J]PA]+0YJeEW_,.5c(JL8[LL@dL.ST
:^_S\cfM>RXUZ@XM>[1.dG3CB,&S9P=4cCFF@f#0MX<;3BU^)/ETFQ;ccZVY\5a5
VVgG4d(;f>NM,OA6+,2+ZDDC1JCEYJ2Zb?eSDHUC(0g?Q@\92K7bD7Z.:3Q47Y07
8.]#89,PUJ+e/e)9e3[f,71NH1E#_YL67OD@)Z&#PFW2O;@Od)9e3KJ#+V&48B8Z
&<0+C#RdWPdFP9DAP@+JHY?#WPBQOTO2>7L2NV=E5A7:B20AT4NB&_.YOI;Z16?H
JW\Y0\-/GQSJ6G::HbOf/6;6fagaZRYWVdSC@\D+?(;_@U\4AKa<<9dP5A-3J-A6
U^JH[b45&9Pf(JKP=]&]/IeAS>QbY7:_W,J]/SQ<Z>L/B#,@N,&)?X[[E\)M^6?T
]3U<]G(Y1N_]DQa>G3=ZKdSGVe,5f(636]SSIfID:GL:g)P+8HN#&eDcfEKI_/O-
]^G^.]Z;DFOAfM)YPbG\-.3.2V(&eb<+f@J8Ag(T,_/^(GdI6eW2K2PJ,_C[0=aY
I5fM6ZAO::V,X,#+f?K5U(R6TeL>^C(WVGN0J_HO]A;TVX/1a,Y_9@I0g)L-4bd3
#0S3MR;4F]QRF.a9>IQ>FLL_=&]1(_;faC((dGdg6+<]0#BI02;aX(O@3_G<@LT=
:CLbH2_IT^<6D6L4#8C;:D[]@7I=.319J_5dN<Y[+7AURFCX)ZADZdE>.CB#7UAG
5D\7BC#__8]RSSBFgIFPeW\e057+0]JJ[(+eQ<A((;S2XA7&_>?]5Q_/e_FEJ:,b
)YL)-RV&=C0;/Z\E-6#RA,EW9\[+AY.1LZ/N+R>9(^8e=&FH8/)]bQE@N\,QL\XL
;6K>V[30638Ib?-bQN&AH9E,6K-RNF7.(aUFDd)WPI0Z5?.f&@7aAJF@L<#O9_2F
EP0L<N^5E,EO/(,gD4cJf6=46d1E.[MVQU1U>a@F-R7MPG&NNG):-22,ET8:J1_H
JB0QUNLEW\?8_EJU^.(U^9U,\(<H@/Z]<N\eIa[^49J?JDbMUQgO/U)EX#WIg?0X
=15+FeJJ-KA142dX@GH0J+O>J4@4<TCb(-^^?Ga:cGIdJ>)_7;WQP3=(YIC\eLN8
X+=4[HC6DU<:2E]b,-WScK\LY3W0NO]4<@B:LTH#2(2&+P;W0VeB9)+c3[ae#VA\
]SPUY4D>B)FR+=SZ.\>/7a)VZHg8Y866(<9SX.c;-JR/3<A/U@R9-6,dCJLQFC/N
+>TT_d\c4#<XcF2aIXCAAf#.@C;KD>^45)GR04HZ;P9>XeKY4gf>e,5JNL\8_a6J
4MM-B4-b[<A>L7AMUZ>;XR],].#8WbRW@?VFPPa)?]bWSG)]:>aKWSRg[QVd@0>/
E/O<--O+d&DSJMALQDENCQTM)B<VVU;53ObId;7?<-FEe1-^WXW;_OIbG1gQIMXI
(7_8A&I:.NN4OM.7_:R->,9c+E,<NKHU(:7a9PdJ-<aGeFFC2Ka^]8A5XS7ReF;T
3cJS16:PU@W]PN_R8BS=HPQ?GD=DQRa/+10,)=P6(9aZ(e&Q1W3MV9g#>-@B)F6;
)e]HP36?cQ1QFW>YF0:W+fXPZA-V@:aNAG>VB-&fSL6L)\R18>L8XND#fQ<EKHgS
[<G]:Y^3@_07b^V0C7>/XZ6R&<.VPZ6MU]@SHDO\T=7/Wa,?WY/89^W@Z342W9VW
E,G@3:NTAE@XDGW\T/-IA9-FMTR.2[<?[(K;DWPTMJ008,AcS4U)N6_@9FH&I?^e
PLC7c)^.T]g),A;f4YY4+F;acgX-@Df^?d,&??T7a>8D;QD45VB<7V&+D&#HX/E>
ZH5BGfY+@6La:9UKHMQRX&[1LeT8\..-3_V0H1c.:<M9KK\Z7X\Q3+@T#O)GBQ:I
FMCVFC#Ybc(^W]Lb/40>G^Z+7>-:_a[P^Lcb+.KaP),:IZH:5T=@<?F:6.7#?><D
T9&,5^I0SF3&GHUZ_OX1La(:^Q[P7G5YI<aA55FXd<FO291c\I83-H(>WVOLTUIb
-R_[2\F,,?R,B\4MNZ6\3f+ZV9U:YHF^/0JR<^:RbfO:ED^:fU[3XQLM3\=MLS@B
0d>VDILUCg.-TZ8T#MZ5b>PHNP8;L+:B>>[EG<HV41Q@GN./A2Y/6;b<0@(N#EbL
\[UYZgZEKE&6g>IM)N2;7YT)^I=\gb:C;^7Q.6XVDb00I6)O)J3@_?X&EWZ-,3S4
ZPS.RL8E^GZ<0WC;b/6(@5RFP#@&aWPEPb7R<NXF/BHAGNNB2IRfGX<KYIB2NSBR
]#c2C,GZBHCL:UH\0XHdQf+?(;]U:HL#8O,&8b8Zb.I8RRI2-:V=KJ7fUeZBHATH
g9Y7S?)PadV/7?#>B=C\733fObN,:-=b8fB_QcHaf4&X^^\b28;59SCC#>dROeS1
XUO8LA,U7VbO&&R+d[9)K@&MHW)B@ff[&&VcKD7SQ[.fSF_9-0Sg(]B81XZeF3H2
@8#:B2J40<5RII[C-=G&Q/Cg^IAQH02)FL1Nd;)6P&MBYW_]^\U-(F:g/bd@gN?_
)C8<;Pf(HI^aaA=2d,[,FgXe\;H\:R?>9fdA));(c^TBI/X<gE[dDcc#S49T29MF
CLe=4^geK+d&99J_f@a5>9fV8_+<8;aT[>8L_f.1+P2@89_//RQKZ>/J<Dc<7GOd
ZdU=+VZQc:e&^,gbA[Z6EDM(?P5I@#eUX43bISM+Xf4(@(44_I9agT:)=I_F];PT
d:^DC,e.G\D/\DC<WYYRIfgSEG@T+;=)Z7:Z?:Xc@b_[a:\_MdUd?EKY2QX/:/.#
WAML/0PC:<eUe&.X=(:)b4c1@+BJ@17g0fX:SNb-Dg9#[<aaE@GPO,aZ7HF#g\SO
dT^0=N0:3ENYXODR[MTdTW)dEJ>@aA+.:22-Lf&&OERX-Q2]dWJ,7I+aH(<BI?9J
UPS<4?ATU#40Q5.5:0cHM>_T1^g7/^D+\[7C[K=XH1,U50\K=,=e[WMW]9XW@_b;
Q:)E/<98J]Pa>Od_b#K=Q&/+NYH#&WFEe=_W>]fFPB)GbA-L&;Pb+dS5a/QIJ1^H
&O#+/?.0cJJgcZ+f\4=.(G.L\g_A?g&7G\8:D^]V(VaeP@9)U6IW8X]MB_F?K<A1
:#TR2&9,-&R-YI+7:\A]A&A4D[ea]H<^X-FgSQ4Z@N2,ITM+7V,UbMR/MdCYQHT:
QZ(.)RW(MJ-e94K)I:<UKJb33dDP;7BGBd157HHJf/]]_g3ZR8O0,5Q0X8dU7;Q.
B<1gB6JQVBgB;XV]\\0(9,]cV2]BH9ZX=@9UO]:(CHb)FN#())I^9Y;PW3D&(:6;
&dV];:OI]\E9De&LU_^(Q&T+1-#2,^N7d+4<RSeS3=e2?0[(Zb/PL<<,(D)<OC+O
WMQ(XE=[=2D&/#cX<0P,FO[a/Geg<)V7BVCeDZ\aNR6:1F5@OaGfWVJ=R4bd6a.M
R\Q\B.YQg1KY/e,U3W1,#CgSI\>+]IM&-?[<;<]1c\LU-O0e7A2A>U-bd8gI[\/G
J0Qg6H58VSJ;I0N5D>AJ\/8a9-a2I&8_H6W#>J-<fP5TQ5>?V+TW2-:FH_=a?aG7
/^E,c:@FDP3MRC[]V/X,Ta\Of8&g8;,N6I&^UQ[1dCQ.&ZPL4g.L:-O7?A,bdO>]
N>C\AS[IX#5]^(3P+CK#DPI_\+K?)J<:\I^_20ME;>YIS8bG\<:,.[CK(@4(g@WD
_^e@BdG_g]aTT[CC5X_EPLP^54K/S5A\EB86O@)]F;#M>W<_2[GC2_?GV7FQ5GU+
39/7YWe0<T,11\DT10,JI1^0<Bb-IR<\/9Z7V?/C113g<TV<1TZFHZMW<7ecd0T4
bdG@]E7M?g1TGcceMHE;fAX8^6;[SUEPQJDddXIeBc&2Cc.-<+596Qb2eY7Fc--8
-[74Tf:VD-GQF_.+G?@PP1M0\Nag5W>+VI@+IKY0c>7M30.[SF0QT+dS./XC-[N@
<&-2+gA=e;LW1WdNc>;/bWIT>(:,+I?E)b.;#Hf-;<,_aH[d7^HOJ2JcY<+WBF(;
1D,cN=17QgT><O3^3UXHM#1WKL?b:8AN\b^&DNN::?J-7T2T3,QR-:E?4bb);:Ub
fSe<\XXEZ73RQYfC;05+KU+#2)Ag\OfN0ET<6IMLGdFSN;AXeY&9:K12^<Na-Y66
M,3a\.-g0DHPH3=-#;(F7)-AO=_=#;/Wf^2cS20?[?UXEX.4?)RR/UZObd__N5.W
JZcUHG]QcHXbJ@1KX^Ga[?RTXG(+_^;Me8@Zg[9;Y^#]3QNAAJ?#[1I;JK1Fd:d\
52F95IDgYK\4?fE]V-QE41I1dYX?BW(HW>=-<&We_P-U]]P9EE2fF>[525cL155)
RZ_?FEV218K(>c[eL7DG>)#@5H:8S(?;gKG_@LN^+BP)W?3)43XG)7eF4</S,Ka)
T[NAT5=f_#fJYgAUId0YWb?#HM1AW7=AS/6>F3W^Y4^Ba^0g\8g?8[[GeKX98-#Z
4fY:#,ZE+QdSXfK3d#Z71<,Z+<81Ig.,:&=Jg^1cFcG:7WYJL?I6P?F,a<<E++XW
S-?QFc8?-+5d3Dc(V^7I<:[E-Z<3fMc\W/1BN4?O<G#:^X1#R\YD?EcN:P@eg,AN
3Y0S>^J1S4)Q[<)ML0^FC/4,:9#).RIaN7EZE#OVGI=X1&N3HT:[,[I&c:cf^aKD
NN#\H28R?QZ;KKA7T01+^T3(^Jf5/)d]W,&EG__<X1OP\-^SM]XUJfca2(:A7+=&
+82#7bXHE_?Nda^=TY<->QcaJ>TQZGPSY4I7U>)P9A3f&-N>acO_)KJ68H@0cT:]
HS,Z47P^(_[OAH\EdR[VOVELF,(=1D^HO,QAWA7?d,ZBYRg/YK/\g5U?fgLbF:]^
R01)GZK^J\43W5_3B-0d^.WE[4TC02@-d,7;+:XTdeE/VJJG<N?-1>SbIQ]Xa88.
6B[YLUd0X>R;g8NcMABFY2^&2WCb:8JVI;G?X>PC6/gZ?NZ&=4fMdGA?O1e+V#W7
aB-<]MW-BUI\bg:A0dFc\FeJ?&RMeXI^ae-/WX9V;,.g&R6J_,-Ib5]Z,UD]O97M
a3Y,8^?F(/6IFd&e_50(:Rg7aF;CW9]HB>9(A3A0T,b7,XU;7M\M1WB4PINe4GNN
QS0TG7Rc8-#6L&7^GS(78<,>DRgfO7YS.bLT[+:7c9<#A)B3cW](FB(+.e7W1Sd=
TBbePXGe.6W__.[>f;?+bMcZH<Z&B]AJ)H91K2Ia)?,6UbMJ_=T]GG]Qe.LF&<2^
1TH(;LeGY5K.W&,784_FGR3fSQ89e&<E5Y(E/H]I+FV)f@gL5H&cE6>MJ+Fb9P@>
;5?5:MZ7M/3-^b)N(^Rd(CXR[&G.:b5-1(CH\8.>;XW8d.)-G))<V3QUdbRM^8VL
7<WWc/UN((Y2Z5Wbd_I[AAZLQFRO\FL^JM(.d5J(AJLS.TQLNN@&11:=?B#@0M.=
?H816V;4a4#BE8[,;:_NK=F7b]LB_[2RR>-LF.E<8Y3,:IUeG.]Te@)E/4=<IN,\
5,BL\T5dTW2+Y;F,K00/eM=,>gXL.9JX;9459FM0MP,KPYM,]:H1KSXg9^1ZID1C
VJK_#G0X01/T8e;--UZ9\.b]V[dK?K91g9D.L-aBQ:#^8<SFC-#+]>?&EY,a;,]2
SN9=8bA6&/6KZ7Ac:c::0RSaeeH,bCOF0;_[XKZ>c<>3\K+=[=D1I.0RP=UgX?V.
RZQ#(g[>aN:b<4M()NE[5b7bSQS1+ce5F>O.&PVI8VdReQVVeR8PgLR7?8A9:F[S
^WWH636ME;ZO<8SR3O@3&<3/B6T^GC?]G3+e6JM8Vgc\KD.Hf[2fY?HJIg&K=T2F
IA?2Zc3D9214cIHf/)5<2Ze9_:;7WN,/>E,_=V(g9J):;e@/=)c=BU;^(WGTX_4E
A?]Q0<&PE>Eg7SGM#T&D4.bL(M^#0]K\F_2e\HP/PF(_]&=;_T4;1Of@fJ)\.XE8
7ZCMC?5=4<cGE>:R=:UAU0<g@\4^?Y&1^>/-fT^73TL/G1BgLc_H3MK_Y+\)T1,V
WRQO6>O216_?>ga48=-S[U(0d^@CZ<N;@7cb(7bFK1ZG&)d=OX>dHW[]1aP,>BRR
:IVI+)GWab\5eca8A=A[^gLU/?F,@Ob\>(GGHRVAH^OK4L3?2Yd_:bgXNB)=,O>K
)[A&fOQ<cQ:_;1JJRBV@aMeU)?ZX5.QbJ44ZO4[NDe0e#9dcM[=_\_N)8a.&4eVX
Hd;:WF[W8[Q<^O@CY0Y/WYF3X+:@S03ET?+[BX48?,EN06NJQ?b]&^:aTO?gA=\X
K3+dD#4:UE&Pa:I[ELE3K\Ig(-feEa42-^NSCA_81=BWARfH=,_E+JAPJRN;0#DK
A@RV1S?gATR<Y@-[\PZWg>7&g.Y51M<T=aNdE0a\^A1J.H&14&A\a5J=F5?,#_XH
GcM_@(8L\,,^G/LH@FZE<;46+bGHV1AdX=QRE8LE@Q-62gdQS92OCZ#IT-NGK7YT
=U88B(42:cAf]cAE:6Z.9Bc;550_WWLg\J&f1TII]657B-+Dg,VV8SM,,0IMNK9J
GV2(68)5Uf38J.\;,Nb1V;g.^[]9_U6D>Ta4KI<47A[(A1a>e#USaS.f,4IH8_V/
Q<<8/C:\P@=f>JXOJE^YZUZCQY2U0]/KCZCM>RL2[B]aX\BLM0UdS5-T/cW)]CDZ
0.V4NOAdF2>5.[@)99OAY.+N<6U<A:UK^#GP7OUZed;(HILUXe1)5Y.6HdJ?f.=Q
:2I1X9dG8R+H91NcSKc=BVY[M49C(fK/5aF5VYd[>S6g2fY6@I0Q/.Wbb)5I^29d
<9gf@(WVR9EDG.L_]/d&c>K>dM9P5>Ra3+(4L\N_@?.0d_,d6)/7C+D-ABDA&N5<
=DGXJZJ4<A6X5NHHJBeK84=V160>6AA,6G?]d[@RX>^?4^.Le?&9UB..\3LC,HQ0
FB4EOG&d\<S0\UAZB;aY8b]]\D9f[gC<YKf;[&:=+[6Y^+Fe.M/-dXfJ0,)#31XK
]]N/D5bDb&4K;:fWKB_Le0\>#Oa\ZVbSYMc/)D<gIM7ZMa4g&DJ@(2TAQe2RCFea
c&RA#/O\Va+&]G>;VWM1CGPW&AM)&)Y/E=(BA^[7[U&9/d8E9?eGK3UM/K7g,.)@
=LI^<\cE#GP)ZFb[D?L\6)eWd8A+HO_QV&FL)#CZcF@d[J-P[VPV:F.C9UMg+2D:
7JUPN/Q^@9B00YY+Mb-Lc;9-QB::-I<F=dSLdEE8??Cc=(]e[YFA>Q+LN=P5K^MY
G<BCX>MP:,G1TSIU<(^HT)]T-,+#970ZL0PMO8JFHOS=7WH0/SXG8C&+E+<;a761
5+e^H@WX=[eOR\?9,351O+UfU)OF8:)\E>bI>HO<W@<2F59V6G5#Z[)4FA#&\?P/
CH<62/R0g08ZCIYT[M.Y>);3]]fGHR?c(2JYfgA>gBd5RAZAc]Y,2-VN5b#4)8Y-
GYefb7A=^+)BKZ>PX(,^EM3MI7H?(R:1+K\^Y)<YVZAa5X6.XCc:A;^7Ic40Hg:J
.WZW_7#R\T[Z577YE+J,f#;=)\U9C4[=f/4)Qa9(#eWegQ3HC#^D#Y#,M07:ZA&(
[];S(),<^DQ#;E]KK(X&\a-X:_4<:?OAbY<DED/C(8;Z@?HW9.]C^^B]Q>@CC<V<
F(=RO[1^:;=YXS\E5,Cd^]bLf?,:f6K@NF=Tf+ZH(cYWX^&R&;XH0V:K/5A#PcbQ
H,(ZC+0,K.OP<-Dc#=-1NX4P923K@-d;1,@?9gg=7CAZSH4aPXQa/^&K6^DdF_],
dT2=27KT_+D1f8F9MZX:FJ#;+8?J&GgQ_DN71-]_cMC/#+g1gPa^-YE&S#\V)MQS
f][P<><)N9@V\J\M[XPKd;Z8=Ac7C^ZCX&&T0X3/&X&K6/[]&+@,\.Cfc@0K5=O7
H9T,IX1B-aTg8U-^\c6->6C+d01HDT3-6?5#ZH8I+7,)RPcJDC@g6<Z:Cec[:K\S
ObU\CH_E=fT3)V+;/3MV/_EKQZ:KN>6U(XAXU@(2@F8gf#]^0J1Ugaf_+<,8<.L6
^aK@REG7&;P/RffS78^A[7Q=>GI081_W<AD<HM8^YCY6CM?9)g&E:Q2gP0XU<]0N
b>JRa<X]QB[aVFHV0927,d.1DJd-7.b;2A#8F,)7G9UYGgE_.G0()5=b<Ge^@^X5
:bZZK5_7H[05@O,faHGEP9e6E;VHG9C8CJ/B;\3[-@=&LOJeOE\);8Z5YR\[5a;[
96W,_3+M;XCJ/)=E8PD/KWS2-Q,7;g.0OAe^(Mb79GF;UZM7,=e,W>J8H12V0(A3
73;Q@645[V#/06=-ZFZd;W)<,bU?BHRA>O9JeXcL5IX@^XK80P_e:FEFXWNT/<QB
MQ]8]=9X59Y>Db68?[Ue&&_EQUF&;).-,37HdL(^TeO(H0<NU6C35MP4,P\-F0]Z
Z7K(]1eNMIgX^Ma,60.6-X)7Q[@a=8ZA(</2FEDJU\RE2HB,&PdK.B,E8>L_82_-
(dG-^B6A>3AT5eQLYf.SgOYR#\>I6(6-K418Y#Pgg?DfR0f.b1E27ZBK4a0\LgX2
Y#c<>H9KBQ^45FFTeZ\+OC:#9Xf:L.X8/Q9ffG]<-5WgWB=XKI+(e^Q;fXf_Hg3e
_PO2)^3-GL_0YARfOKZVG&+:IYY13.Ga-840BF4(@eb5@7CD#=TD66OE_4MLd+_#
U^1RF[[T]L44cBG8C&4PQH:eCWc7?Y[LGU<&_Ed0Q)GIRV,RAFMPA7JYPD>PIgDT
[-J<cTM>S3e6\IAL_5)ffF:ebNDg7-/9A4G\2c@c@]cH[e4124E0(;9O)9S=Qe<B
8^[0]G>-2fQ/--8N(G0(4P5[2/_P)dWL)V:T-aE<U6<=g=]&_QH>=_+-e7daF</1
I,T19HN3S-PV1)0H(6FQTL/MZ,K\8140LHY>Q][U3\<Fd?>3Y1KY=:7+R\H>S=(N
I#;JULF1>3Q8ODK7c:)DW2c]R,]U4HK+@R?HGF^IK/[b,=/+NJ_gZKf>6UI?1RU=
c1f?#([5WQXbe2+/VI-9[P94R-9>I/KQ3+c:7VZV;ZOa3g4]S,b-bdJ4FF0>^9;:
aX3O]C58Zg,38#PKd^1>Jg-_H68M^0G<JAf1c@f^cIC.g<YH(dYU4RJNBR7Dg&e)
M:>V\U<Y0:c[C^^R>L/LIP+J.0>eKXVE[8YL(50.P+_BLM:Z0-b^88^/CC)Td&LL
A7Ie;aW4e(?RJ&&aM30&,L_GQ^SO+YJ6AVPWfGaY11:?/L[^f[18;ffeD6f#&[.#
S71E498@HOCP:W(CgWM?M8_PPB6O#;]69?I.daeY1)^22:7&&0a5Hd?5H&+]3-(6
XP7)W<G(W[+[b6BEPK;fe7)8P:L@GYS4)Q+?U6CQc@6]G.7LH7)a5R?0aM,<]]K6
/CQ#3(>E.f0_C:g40g9WUE1.P@g1IG0R9L(DR)NQRS@C1-ENF0TVM5-ASK0P<EKV
B1Y#BWHVMRUaE?VU8\b-82&CJg[:5M]fV=IdAX[WS>&DEK=91A(HH6V4D_L)?N0L
1]@&J?O8NL;;a>bMTdRZ077D\9;[EeTgF=NL;UK>K/@[C+g#\-1J>b+\[KVMLTA^
1QZa/;,\.1F0T8OOIG&V&AB8Ig:dNW:<._AbQ4]17f-_45YIJTK8I+L(=PC/4,&<
.1X[N_b_?a\L_52SgZ_L/9APbA7XbMTf(,dW,@.H>CCK_)?00S@6fE:>:#QJ)[24
P&[bYR01bNe0e8I[XO1@BY0>g]fd98=-Z&Hg8f#HD?Ee>-\=1M@H)]cFc:WUf,Z6
YWK>;EbW)L=Z\SQ7L;S2-)B6B(]E:bSZ<+7(VXZM(J[c15W88RFNd3)#d>D)>S&S
Y3<:+82N#dc4^J?4JTYI]a4:?Rc4-A4_N;,db(2(H).N[#NXYP6Y@,>WJTTaD(bF
U)6TG9g)DO>4JT+?d8<g7PS.YQZ#J<K=<K<=]eT-@cf;4&@UWcaUSKUfKN\<VPR(
X<e3:(bVg4]^RKHQ]E],8?(2g_L[.[(V;Z@O:(V+3)RF[JeQ#B]F]OaIT3L)HPfC
=>^2B[:&0g)[JE],&#=7W355+LEV)7.TKS^eEV165+5I?a[bHF6YWL[2:^38aI\.
W]V?FNZ:/&B#,1<IAJ(g_2+N[1N/d2\-1>b-WD@A#)8ZUUGVP3KKf6)M/5_b)(S[
[&6a:LfDaV1)<Z?8aQ2<5S:U-d(8K-G9WYX/]R888c6,W-8=,&a]:>4d_a<U38W<
\2I\T5-Z.FNf8Pgb=gOXd3dbKZV6BeN60PJ;<3gV;L?POQH=X.a,f=fKIN#)A.ID
.bU6aAF?ZXKH\P21RT49NM8e-)DYHg3SP2R/TZ(?LbX((AT/Pc\_Sd006e(8C5Xd
2<?W2M:\c0SZ/A6[-S,-\T=XIPJcIB^eK=[3J3=2aE=8/:Fd2@_^A^S22\;BS\ZO
6(17LR+DB.4aXUcS5cX]X5LQRfUb&4aT1BTQa^U?bK2[I#=dU4._,_@LE,CE]g7M
;P61/-C(\_I8,J\O42C?eE::=^[WMIL4VMOWcWI7JQQPHU<7/\U=c?UHL&U8\8>B
(Kd14c3d=eB@+WQ4R@_N\LH@c&HNHJ[9L4RWH4OM8?(5SFY@,f-6#,S0R8UQ+?U>
/f4^2JX&b)[7\<UbUL)7WdJ;@E_X0[#0KET2=A>+RYU/-R](b)D7D98Cgb\P;^FZ
8b-;=2L86:BVg6=U0LQR#bK+_Ba_=6/)<Q=Y<F)Y.UB)^_dJ?P[<NJdB)IL;UTA+
I,eR&7fXTOS:V^YF@0(]ZWg1cNY[-0<05:,&e+)/O>^/R;?KI?FRK<FJQ/9<K8Ra
H:#4a^B]:]=(PMWdQ>,LfJJ\.2/CPg6:+=a6Y.?BO@3+Q(LR[:/^88ZJDe]4Y^#F
9Z,?M7,JF;>@K[1CR@39/E&FafdD=,O-9#4VF[IFeR#GIS(B=ORV&cTR04DC-+F#
ZWGT3aDfbYdc42,=GOd2S6-LY805HcTRO,I#efQXZd4B3G<]P+82]RU]5fO@GMFg
O8?3]?Q.U,-aV8.f[9bZeF>SaB=RaaBNIP]9QIgQ)bQWB]6ULFeaS_Z^/#D)7)&0
Lg4B[[O</[Z?.N=WGKPH1gQR\D#GI9K@f;8Nf/<B<Ae;C)R>O3b9X#V_(]RPg_2Q
1\Q=U2BUeaQ-^R-^7WP_N2)+2^T_]7;4D5+cZgRb[B(d7^PeS90.UC&4GZ,+5ZJ0
f;U9dg;Tac8GHAAP8I/@I&ES4/HJ(Qed[EYaCQ6g;cDeA&6/2Rc<PF\\..-?O?D9
B@a:cPDS<:YJJDc\>P]+X)@WSJDD.A(d1M]>G7Z]LJI+<;?&EEJEbVV3-D]@^2K=
DdFa#Ub,7X&1XTF/(+,),78)cX(/8DK[.=DU:<L8ec-N:4G88OY:\H>++)d>DN]/
R8+U-WWK+4_N^a0;?ZALL0&eg^K4:TQ/PTP/>(7=Vb:PYMF(BfR=f\X4Q\U[dFU>
[R)?TNW8M9PC?d3R83@.P#c0RW.:LMa;)]Y/X;#LF6S&(b]=SD.eO[PZHc)<)M)/
JJ(Vd:LL<1HBY^OYfV/W-<H\A9:R8=#M7aE3>0H0#?#/dGMPD<1(3K=C,S.WR@Q\
;5R:YO^X?P[E.H,T1c&+2L2V,7D5K5dgI&;JDPAY7BXYGPB7;f#FD#)_MHIF@V&U
BBf0&Q?&,;WAEa]5/9>ZJ-.e[,LYTAIM^WJag&fa3)WVKc[[[cNYNACfAc8dOT:+
L,VUHBa[F-C0XF\D9IgLOAYgI=-:\37b3fT_93.#NTD-F\QBH[C&PSg&B>Ng,4)5
YKC319\[;=EP^1N)PGB8c+C3-(a@G_)V]0c]5eSL(1MY2b]8/g-=</P0J[,WL]@=
?;=][>&ZH9aBA3T6^SJQd=LgIQLb9<;dF@ZdB4XV\T4fTH.EdX6P]_K]0GWDVdA4
GR97aNIbd420B4CTOZgEA+;.>>6G:@4J9^HE4AVZS.Tf;AXN;,QNG)_)ZbL5KL^4
5/2b)3N>1:FQK&_8g8WUEW9P_C:HBDBEf;M__(ORSEJ<.B6PSH?g3DH^;-2S=<+=
Q.;4JLGG0KSH7KY>1LB,(65T#8I2QN;---5.)aR\U8.]29;A,MaM=X00@XS]gFME
XW?EdOC?<f<;Q5Pd46Q0,bVWabOQ0]a+3X5>86]7bCP8XcUZZX?_2d-E+1&J/gS2
:<R#)BMJ?MaAQBLF1LJ:WK8SCR:Z7]].IS4,;I:H_##1I^3gN^P1R>2\bT(eZ)+.
0c<4BD]O0?&,MR2P@JK(+/RT\K#^bHO&&4YR,(>=I+.;<L<f#I?#1UEL0CGN^Z:U
LU/JC2BabV>)>MT-T.JcUOE9^SQK[\e9TJ:d?T>_K3<^BK#R0_OW32@/JU]d4YK4
-YYURJOd#7VCWZed>HOS>U.^R6g-Sb\:T)#[c)Pb.R8TSM9fTG9;(:#fRXY&H=Ec
0LLY77Q?XbcUO_9R#)P7^aR_)NVa[+^A<<YH=X;HXZg.f@Q,6CO_>e;[AWDaO4=+
)U<W4YG:?M\XW44(;b?1&5+L?C);b:9WKK.&QW;P)HC7]EG6W[\)=T(H6XaQ6B<8
\-NcZIF>\,bc5-^g-J/&^GbA.c,IU-C[NUQZ6#@9(E\2Yc+EX5,B=P@Ra6)<DS[M
)gGRF5c[;V6A6:(AL@0CE(-0H;-FD(cY2QZ#^3E3L6dR#\^K+=;BS>)4-2/_3MM7
+DI(2Q/VbU-3V:^E:eb^WdfBG;6Y-+-KBJ2A7#J&D\WI@e?7:HPS0A#IQRXF?\#c
^XgcN^.)^E7a@<,0e14L3^8@??eRZ6dLU9M\aQA6TETX>U/C1Hb)e+-e)0VD40XL
;HB,Kd.//M//]4XE]I(+AYIQddgN?^_RTJ90ged7NCDH#g[[CULcDC8S+8E#VT=;
9I=Z8(cG/,b4eC#/bZdH[D9Ka;K[Q86P4=cB\.3U&:R5@PB+8PMZ)dVSPULL>N2g
B02;##U9=eRe5_ZL=,?Mg:e;9+MGL0\Be()2W@=H[f/<UdKg@&\I+MNI186.B;a/
M.)Aed,/a(6E.DEVbL>e=?EegUNQaHPF0.VgP<PSf@L6-O2Z/+K7#UXV15NVc#(#
]Db&33WX5--Pa^XD?QIgJLe?Z0gY6B&KXUSFJ__345O0B@88S)H#]gCBfN8-d,#<
QBN>^,^Yf<V9Q^=bM]_JBE^V+C46O-/EQOgYK)ED?_U6(f/X;:6PbOcX3Zb,5TB>
SbR(Q:5PYM:g&^#IN/<#=dFDLC8EbVUg\0[cb(fV?-YbFD4cJ]T?2;BVC;.9:#)4
_TbK94WURa03#d.[KL9(B_(>?HKT?Y6K#5T/JIHYA.EUSDX-)/VQNEB.^Xc;VUa:
a1ge)4?b^6)QI;;\Z=5/8YA45ZRR-?TA9&]E[)XMZNeQb6>D.HcL>1B..Ya1R@c;
[#:.]8?UePUDT^/c;LWB.cdZDMFLU>>A4fbTWZQ;M<-<\K[WAAFd#K:#_gEHYc3>
.;QK\Ff?WD&\H^211aG]KLB_H>a\;RB0+J,LJIW[&2-1JESX]=XaHc1_P:&.U?YO
a3?6-436/)6)0]Va?=Z&3038^PAE5]BFbM[dNYG_R>]:FC[56F-::D2NV])f;+^7
X-1YL8.=f[d>E=N9\[N<V,VFVM<c;=-OZRH:M\K6LcT7V^6=e-g9(a,=5QQ:dBM]
FNGOCIKSbM6D:Z7#LXCM1M#fMXbfX[JPHbX/#=W)U(HJ77^]VH\;M#Nc[1Rc;>-N
]#E/WPP:(M^[U^W@1J/8G.<C@,f-]GVEdc[>A.g7c;/0Je7g(/aT8fX_A<>(<-Q&
,Uc@(B/99AB68=#+a7)NA/O92#L]3O-ZVRC-TO;M9JE<d9J^,,F#?Z&[7@A42)c\
DP1+gBD[-&IWRY37SbdYK@?2e@bN^\cQK>62C>Y1dbDJ1(Z+Y^IW+Qa96#OP_PdR
+]YPD0e2U:/EK.,Y=8N@a#[AG#I[J+;b@0WMCg,FU0Ef@Q9X?A@e#KTaP1g8_F.:
^U^]NB-dBKA^<7bN2(QT#&U<C?03gMXFG@PWSK2&&7^6Af5J6DD>?D5+,&b)+&_6
IF#\;+]ZVLIOVN/O<X<.MW)fX#]3BE8G\g(b_Z,dEb^_7E9ED-4S5;K1_I80Kd-N
Q4;6gdA31e2>Zb/acO-,2=a;90TYN4L4QILC8KMf[9(8]WIVS]<K;WT.88b\N]b1
Z0O4?\-DfHY\:DRFWgI_YAW4)V[G^DMAG]#^EG)=Vb0SX5Ba6=ee5T@2P#9(-1C>
]c/>PUC&G.80[W?0L?&(L>N_=T5Q7VcUB?5BFLC^BN:<GU8OLM]d@SOK3LG62UBC
MCIC<U/TH13UcW4D4&X_W.La(P_)64Y<UD=aGC4C/C260E89QDRL(MZ+MA@(Wa;C
P<E_.7+,Oc()<9CM2D\I7,b1<]5)\1F2X4JXEGU1.GJ;(AVdJAcgIL:GdS47A>4c
ST1(U&^+5M@V=H_\VYO[9.M6gb^AS?C5Cd9_XX//E^EEN1M-Og],g<7bA4)\#KMJ
Z9,fSJe^(/9U_,P[0D[:1Y_<>g=D0TNO.9_Ne4I2?IYgKATYBf>+O=C^ObafXO-G
6QDYJ\\WQI,GFCMWY;9/:dQ-9#RUUJa2O=<K;9XKR8>M[XR@eD_3AJ7@NJP(_RNI
A66[Z_b74g?-6X_?M^QR]CdbcK15OGDH3d:.gW+F05NTGg-2e-DG]#)@FJJP?H18
.P5.TbI8RYA\R-aedIT@YNee;@))#,6Mb=G-RXTD&8?c)FEJgL/dAO3F9UKa^fXR
8K^<3@fZ00cG//V3-#P.f2^8/EA23#QOX]&LN6F1<WUdD8C4SDU#MHX;2Q?fD04E
@360L#AHY&XO[<0ZT+RUW\[J].IPY66fXb9+@bD2>OBXfDaF:U/<=#(Wd&b?A9eJ
[F&+JMggQ\O<6/2Q:.R+1H@O,NNb+[,Z5?Fb7/:SRAM=ZGT2=<R&1,<V4M5R_PcQ
fb)a0T;==J)]3V-GP;5fY^c&,,gM0RANB_3?ZT5PaZ=O63Q8.,J@:P75LF0IDa;\
a6JNcJa2F9)&9X95e>QF90@6bMVSD8[:)KAdJg^JWge.aIg6e)3V5^K^N]Kg?NfD
28SK3WfKJbMZH[fBc>c_6[Ubd(5#HY[_&>I(#@N=MVAWR1,N2A8/gg)d0E2OKG4]
E-L/;\+X.a9[28.Q(=DRRD<Sa8KQ,6OXRKNBZC=bU9W66D[L\I)RaeT[+-C/[4Yb
HfPV<WgXg0Y1N2;+AMaUV.6)VYc[A_M<CVfc@6:P=b;MP?Y3FI5_HK,5gIFd4946
^UcDg]2RS2E?85]W8=-7C?1@:XH);.U/MPQZ8.3E_((X7VWaUg70Z;^3c&+^QUI<
/RMM&#/Ce+;N@8Q(59_Y]F.da:K(L[>JN52;CQM=C[BY6(Y^dDMWf(ADG[/:JS\(
3IE+D-NMOMB.C9c-ca)U^6#GB1PbSg7,W_>c<+5VZG:93GH]&QEA1Wb\cUSZ#71.
_Y,>egXI,0X]eOX@N8>?Gg+8b-5=XK<DMeF8BMW3gJ:cB>d\PCNVYg-&YbG^dNOg
8_.9OI.Rc>OV+f\dXZBaY?QB@0L.5LHY-6bKdGG?K.A98OO6PU>?cX4T<PG<1bQC
A?-dM0U]2g-P@:KC#86^Xd,@LYYB=)]gR;ETN_&^2L,=OC+0NCX(3aWSHdN.M.4#
eXCX,Kc2XJ8Db.O=LXBN8\=Cd-<V;MR-ZcFb_M#7#3Qc4KT:A:,WYE(YbRUbg8I7
KCb0_T#3JM[4,&>fG,;Zd/HT2HF@446V>.WKb39_Z3S,V_WYcMS\HWIQJ_G.:.4I
(XOCVP2WW0b0DF5F/4F-J/8P950#e(G,#ZFgJ1edAB.-]O?K=:<S;]aYEdTJ#:1X
3B^CNaL?DC?/D:>-SW)JRZM,fU&Tg9F-;#@&b-&NXRHQ2R@GMCV>^?4:BE_@;f8b
\GMfGM/[Y2]9U0fYO3@HLSW7Y9RJGM>PA0EZ:Kd>?M/cdW-RV4(2G=8VEKFJg_]/
F2YaB-b:_9WNf@+(aSQ\[LP6a&QX6NKG:+.JaU)YQ[:\K4.g[DPCZDDJ]>AfEN?&
M647+I)VC]\<d3,UbQd0[dJIdDJ?>a.-ZD2(CYMX@NRI;S]DUQf-,N^f<U9YcP4L
bW)6@WF5\/V5P620>f\1&ZJ6Qg]X?O7X,>c3_ST(;/T0Y(Q:c&WUTJ,6:[[Ee&MJ
HGcF#Z-eV1MFMf_&KWJ/<P9##d<3AKKd=MW[dE0FZY61K2,9772\BMAA:.f@)I\1
eUS\6<gV#aUVMBZYTcQT_d#c)H1U0/f-UR0QJGPD?_73g4]HMD+BUK1K1aSbe1Eb
g/]R1Dg^?S3TCN;_a0:L&CJJdc7L\PaD7aUc(5+cT@I;MGW==/f749b-ZVcUa29)
,Q:+^:.9J6?#4.2(BETW?6&dXXZ<SX=ae5Z)ScWQJ;OAKV5ASJKN<gE-LW[6A)11
TWVQE9MN#,63eI-&::^K)]KI19_Z(6H3-6FAeJ?O08c5UH5cg<^71Nf;-dKIRMX\
3:E@0KM)@J=_68>4b/EXY&-X1G=SGFO^KLI99\g7)==BCSg>5?f0?V9[/LQWA<]G
gcOGgK=29[7WFc53dC7\.3\[c22:^)M/DO8@Z]gD#?<UaT5gIM)N)B?176f(C#(_
g.,Kc&9f4Q(4G#C;E@TcOH9/g<MAB([c+NOQL,7V6gF@2X1^2TOf=GIAR[).1IW_
W9,364>a7I>^X[AFL2D_K^6dX)agg\?^L4-JbJL6d?[,)b<f4b)MA)TTc+4:YGH4
>90-f8:G-LV+9,MX>491GW1PCR9=E@Q0UK,J.T0GbB2HBL-5FKE;P+:bEPRB6bD2
<Y_3OdZ[<T-e.;BU@b,Q583a<,M+?T0#XSQfFD#YRZ:-C7OOUKYgM425K+,C?M?L
+CV+KJbFV<HVY7I8WK6bMdg(^9^63Q:bZ[0TAZ(F?TUQDA6]e5-Qfe595);WQ7/Y
49c1.Q.U@K.>T.39.Ga]LIRIc#=/IBS0gID\TKK,(-S^dIfGOWJ+846+X2;J#ScS
3R4BY?HK763+.0dJLO2d8ECHg(+T0,T<0_5<e<Jg:,P?;E)8bACEcQ4#83DRLHg>
cHU?dR7T-P).LA?0QUA=df,Y#D>dF6M[IS1H(@2YOF&&LXH9MI#WH]+D,]3=#gEO
0.+H>R,J.V]fd:A=^VbdXd1H<Z)57,<MeeU?#)MeRK0[_SbYXX6(SF3_JJ+-7bdc
6/3@8ed>1BT=^f--A)7VTYg)b\@KOL2(=?J9deWMFcbO)#@GN]A@N5LF<\dR/PMK
5f9\GRc+H^6SA.8I5gY]L_\YDJTDX?C8=E:Z)\I.E1#=BeQd&I)2B<eZe=4UO94b
:&dS+W7]A[eQ-I;5][JHJa]2I\_/RR=\S?5eKgKB:ZREg@L:@dMgIX0]E0^8E>IJ
6A-<XF9:;WW0<I?&WZPA#4C]5O_>.7NQL?cJ(RZ#4[e?+7R6DIXLBgW-__58e>[[
@NBgA@+\0QLZZYfFWA5<F6LNJVd#.3H0-b82>9c3(W?Q)Q@.c2HQ^-?P(dO;Ha3/
QYCcGU(.c/H#=)&@<CN;Zf5V],AeDf)9GS3[\Z0c),Z1J=8FbYc)c28Y@fUF@/-<
US5RMQ=DgJUW1LJ;Q0N/f9H9FO069;ZY-KF<eKT\3\8KMEeUVaYPbdQ#eM-LCcVK
a9g23OH[KSa)N]?1(d+GUM>#dHS6Fg^aa#U(C;-LZ:0?\ceAK<G/ZVJFKI3Y,J7=
IP7QN_6g:.cgZaI)eR.G&&V3/84B0<8RMIB5R=:V7^OSf,N>7b(OV)T6FMQ)b@Q\
;_+__SL7GB9&]/ZgH?b_0B[55QK^_X.LM)F4bgd?/;O)D5b8,.W6b)_4@W&E[^Md
?_OOF6]O0.CI/Q3R3L&W[0IR#<da)RCUH.V;=ZAPT7Y;K>B^<JDS8=7,cfVWNg+H
02c]A^&FaZgW#9-ICdW]ST?#J98>cNgf[Zc2F8I@BNbJA&Vb_AL5AQEU^F]99VJO
947,^GTT+f(=B<)-:J6H<@dRLc8>aGG+.c:1U<MDab:M3U_5^+IWCOBB[S8[))_C
5[8XR\BRZgBZ>g[TI(gG7CP/T>,5[e1;ggZZ.QdgOe.bIV8^NSF:D]_ABb((WC(E
2.KRANB+UBQa:9>6[aX]P353ZA;&#K\N,@g3-Z5.-=S07Ba8)&]T+[QUE3^&#dJ-
H96-7AR66[YB^Pad_^V&Ub_0/=0?LM4&[S]A:H/a]CPQSb=_.S9-9?Z&/4V2AT?;
Z9QG#/6,/&C?R>G+X=d12YE&MZ>YV^)>:RV7=cERZD)EVgeN/]BB:g4G@BTe;BZ;
1E:8TeSOOS>I^&EU@aYI?W:U?:_#Kb/KG@LU5YJEQA/3,@+fc@BJ7Yg)\S:DCFA+
AR&KSg;\b_<WbAL9eXDbOFX]/:I@e2?@A.ZA0ZK^Xe/R14H^Gc;-W3g-+8+3WL,_
B1=6^5.(I37H^&VP&C^4)LVOZ6#;YdFV]\b0QI2eBe&Z.[TX;\c.L\@DQ9U-4]eR
dDMVF);FRD=RLU.W-(KLFc:QgRg==6[W3C)_;PA9aVF(T2Jb+2UN5aCPX.Y,809&
a&Wf\<A0JD(P.gXA_@]DNE5VA.D;ZH(,--JT0MId<)MAL<cR?T7(9#QI:W:>I2RT
-3Q]P)M[6:LN<ABb@BRH4g2SQB&(df4<:aT:4&US3:_NIZ@,E;BS;M38CNY]G&Za
I6d2EV@+(>4Ec9\.IL37dUY)+3)?@Q\-DBCD9WCA-U5Sc/X91S6=)(T2cW@H:>f.
NZ5K#^ec]e314X#gNXGGc9MgPId+GQJ7(]E#B6J3Jb-b6-K..OGU4@\M&).FaB_?
aL#+8L/Q2S9b:#2B)R=3;+WIEU\eV0&14^fV[YHCA2N[-f(,VZ^,.9T&I2c^BJFg
^S)08,I,Y&ec:&0^=QgN@.;b;CQA9M9aIOIaeFR-8E4U>VG/HWd3W?&g\Z,d->N2
e@1;=+f&S7F&?fAG(I?6J)Ag]D+0,4/H_-R_P2(FPd2NKF(@Y_>18QXTbTOPW6PF
Nc(&77/b=X0D3]1^d/dF\>WfYXeTXA)5M7FT1NLZL@eS)1Dca>8aFB+1CF7.TW6=
//),:dS+2d8[;H>;L[&X1T<TXB@\TN6K\)bH?Z=#)TW(N2P/.MPW3H[fYEF].:6P
OUFBLKNR9@5>bb67ZaXH4E/[MdX8?I;GRF])9?K>82;E+W6XDZ2ObC/=+A&+-LUQ
L;eZA:ZaN;ZX@2I-I3-LUfJ&[AH+K)C>-])3OY/^[>ee7H&NQ_+:YGZ@a72)]\;&
]37a&UIgF6AJ^NOb49gQ/QNOV>8ASO=e28)1R)^,\G_Ng3XUZ^^aCdZEb+ZWg+PJ
8#?HILc8G&,H(L+?;E_c1BM:;6JPQ.3-JH3F5H=C/@.H[?:U1,AS)ANg5&c,U9Z@
A]M;1VE-R>6:BR]cWY@c<9@^-db5U\VUG[F[SL15P^>a6I&fE((0RGF&cA:DF]D.
844E/YP/L]4Q[;D.#0gE,a.A=_A3Y,+f+]/_]6<2ZF=#EXeI+Dcf:8F_9@3Lg;aK
WRJ[:<9\T=AVE[JNN&]]9c7-;&aWIIZL@W@:LgNROECS]>0da+^E;A2P9]g;1<[>
^ERL2#8IPYe_A8=)8bF2cC_8Ea/?>.]PP3/.GVS.HGPN8)RB.LC7@JAKSA4J\^b>
gZ[:A(D.M6L_SIZ&:O4X#P8eRL)3MO;F10NI7;03FcA^-?fgLCXH-/U=F&eMYX#B
\+g>eG62#Fe5;?ea_1&gX9&#3#ae&+cXI>(SY?LJ11(,b7PVd3\+1YZ7?9cIBH^C
L]<[WdH/BTW>a8)/+4L-\I&f2_LW[&<6cf/aLaP/b]^f0E]2#@[e2OO79FcM\#>P
X+B\5>GBE<S#6QGcQ,U)T>)N&-a:^2C>A88N:<N\;=-TE?HD[JV3G\4[^G9##UMC
]E,5L]0<JZgeR)FV2P:7AM_@a>gJ/SIJcfG[)PM)f+V._fBe4-?FX>S_4bgeD,__
X:M7QG&egAf7Z0._.BMA7HG<PPGU;ZIQJ+^YD9P@?&[+P./^&IaO#eYZ79Q)][B2
1>S1dG?IURBA,;bU#Tb:>:b.0(7A8&W,d\BT>O[V8T\]Y]<O(fK(8SSe)f=XW2BZ
>--GLeM_V=Ia]]XZ;KVSe;[#IIAeM65LgdO@7Qf<LcX/8Z68D4&_SHS9ga@1@7a]
&^1?L:T0/7eON]_1HS#8&KHFB::>eZ@LS;,E_fTGI]9V=Db?N]D+b>SPb[0Wgc/K
;>4VU4SI4&4RX2<CMRS[QRJ:E>A]J7U=S=6T[32fC0S3&)Ya;@Jg60-&U7<3,PZF
T@1e+Q&0.P6LPRZ8\C&eK665=S0FKZ+BR[,TFgD2+TKABKL<W4?_.gJX<F27S6>.
4RH&=QVLXagYb6dQI@(eZ\eTV.U[ddL-KS#G=d]/AXc0GK3<^S4ZBNZgfdPc:<,G
+9[8#QLH[6(TMJ=3,g3cT-\Gf)a16&9&I@/YR4?0?g7)@#9(]0)UfO=^:-);6_GB
9=7Ge+<RERd<)]+_^ZF:L-_&[Q_;J=()QT,4gb]Sg7FcN2[^?@bAQ7EfaE2?<e\C
gCdMg);MKe+IgX]?RI29:C^N;Hc1BNEUABWJ,XXZ3eKDPFeI9-cN)F2DfLHD.afc
G+DTFZD[YG9T/>/X]e+QcL/5+/<c=fbcWD@/H?BV@9;V0eU<)3G\D7XeN/8ZB@;2
NSZYX.b2>+A27d[fdJa[gQ_f9Aa0)+,fY)_.7R7:A<ad\a^g+AMJ[SFH8F?d<TKZ
a52T&Zgb;c^9M//d<(,59GG5d]+<>8)Q>-<Qba@GWP-QLPY7=A.B4D,;UF/LBTU^
VKb2,CNM#S9XT+LE0I5?gS1,UC#XLb\G-fMK]#E@)I)(WcFCfBQ4D8;,>]0<._>1
6a.QCZ4#_YR5ON=c-X_T):1GYW2f)YV29$
`endprotected
endmodule