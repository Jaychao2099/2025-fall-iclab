`ifdef FUNC
`define LAT_MAX 20
`define LAT_MIN 1
`endif
`ifdef PERF
`define LAT_MAX 500
`define LAT_MIN 300
`endif

module pseudo_DRAM_inst#(parameter ID_WIDTH=4, ADDR_WIDTH=32, DATA_WIDTH=16, BURST_LEN=7) (
// Glbal Signal
  	  input clk,
  	  input rst_n,
// slave interface 
      // axi write address channel 
      // src master
      input wire [ID_WIDTH-1:0]     awid_s_inf,
      input wire [ADDR_WIDTH-1:0] awaddr_s_inf,
      input wire [2:0]            awsize_s_inf,
      input wire [1:0]           awburst_s_inf,
      input wire [BURST_LEN-1:0]   awlen_s_inf,
      input wire                 awvalid_s_inf,
      // src slave
      output reg                 awready_s_inf,
      // -----------------------------
   
      // axi write data channel 
      // src master
      input wire [DATA_WIDTH-1:0]  wdata_s_inf,
      input wire                   wlast_s_inf,
      input wire                  wvalid_s_inf,
      // src slave
      output reg                  wready_s_inf,
   
      // axi write response channel 
      // src slave
      output reg  [ID_WIDTH-1:0]     bid_s_inf,
      output reg  [1:0]            bresp_s_inf,
      output reg                  bvalid_s_inf,
      // src master 
      input wire                  bready_s_inf,
      // -----------------------------
   
      // axi read address channel 
      // src master
      input wire [ID_WIDTH-1:0]     arid_s_inf,
      input wire [ADDR_WIDTH-1:0] araddr_s_inf,
      input wire [BURST_LEN-1:0]   arlen_s_inf,
      input wire [2:0]            arsize_s_inf,
      input wire [1:0]           arburst_s_inf,
      input wire                 arvalid_s_inf,
      // src slave
      output reg                 arready_s_inf,
      // -----------------------------
   
      // axi read data channel 
      // slave
      output reg [ID_WIDTH-1:0]      rid_s_inf,
      output reg [DATA_WIDTH-1:0]  rdata_s_inf,
      output reg [1:0]             rresp_s_inf,
      output reg                   rlast_s_inf,
      output reg                  rvalid_s_inf,
      // master
      input wire                  rready_s_inf
      // -----------------------------
);

`protected
@.;)+8dcD;R-:FO]1@^5e^Q874MJQfGK3-SgeW]>eV>F,FV-WT:f2)ZO-M2E_X(-
FS#\SJHJb(a=9ZEN9a2?AOP],#:f(bA8&Me2JKTD9/EGO3U^\.A78)K:c[g<=gT;
YAR?(GQ6eY1\MLZH[N&C=GWMA7H?MJQeINf0:L,Z:OV6Ad7<Q+RJRd?XK2A?NELI
Ngg0EB4BO-R[;;WE[5)aD+0bgZGfRTJ(&YNAe.>b9[Zd;<3GFJ^:bee]64<(8a\3
Q<-a];0CC/9.f-K=XC+N?WI:U/]GQHdH0Ye2;<5=7ZI-VeQO5/=VX\QA0VV=N.I(
[/PdYNc&59[aK34&Sd\L)PN_<L3S@MZ@(8>cOR^d#:1Ggd2GAD-aE+@M8d\C;)1Y
\5LY2=),?gJ?EWT?9e+8T5XLSJZ;152:KK&.WgIXfbeFIH[WQ#>(9FYM[<d0XM8F
9F:K3X)E3(57PEACGMOeQQ)03J(V[,6U]3=6MQHdV>T,6SgEC6=GEVV]&PN?1_#(
[)dB>-M3Q4G3a64V;,-Z(&VU81Ed(c4R]CZMS>\B:8C@I_L]Uf_G6V,\DK0YgI_0
=0)Re850Zd<.:cN[4](Paf-VI15c@--Ad.9Q>Ag2;-<<(,XJ\([RfL/J<XFIIC=G
.:WNEFX7\8-b/16MQdIUeG=ORN;F:WCDc,WMS6VgA-4SB?(AIM@ZM9COA&I6^\aa
2^_)/N<>@77=6W#+3gH=(V>BAM^E\/,NgJg=d>CC^eb#]e^-.#D(J(TZC]:1dba[
6D<e:=e?X@Q2D/N8(E@55<X/0072D<1I[3(@<]8.-9F70>eV4K;(fO<<37./>J&E
IQ]5daF3XQDYPI<C,R#IQ,aOgGGOFKG.BeF7^gHI9e.B4&LWA.N<aU(R3AKcgQB<
O\;GTC9JGTeSBCQTOBLV:-I/R<dP2X<O_d_O2fC>Sf>3HFQ,1V&CGZ5VKNGE/4MG
2ESc>CJ7MJ#]Jcb1AGB&C^S.C2]W/XTL6U:cB]-[VDgHb/372e0GX/4&G1ZXW5a<
,#,1Z,VR2<f6^Yb:^e#+;Cg3(P8L:;SJDAPfJIS=9cOEJ74CAdZ=6WdT^>-C=HSM
.gM;U8C0BSJTN@VUZ-(8f1<=d/)+Q&(&[?d>3I4f@Te/CS;g;f^13f;;TLB1JdLJ
aXa/Y:dc=+B-K&HWcD3FV0=FLT,BVO-<Le#&1,)3-=,3+W;;[VeY@D;A/+6WcIfG
UUc9:#&@IAGG,_FbKZ&GUE[0)A2<HD@U+2=9.+>8W62UI^A#F\<>ggN@IDDB7G7L
ZYUL)RWSX=6X?7MTGGXZRT/4V9FNRe;(DA\LKZOD;H@a8:AfPa9d:-HHa,LZYC4N
]A0,TF0:)XC]H_22</c=\TXT^]]J&R3<7^.J>Dg5-=U-+:D45ZC0gRI>^@3]+RfT
LUf8_B>K?6JLD[JB/-+JD97[A[LF1KO37c,Y<L8\,.FR3Rfbgf[?LKA)a+8Z7+WH
&/bdKfZYNC^O3PF:.:Z:.,[_-&95C;A7O[IRad0eJdg@.^4d1dRH/0PF@:1_DY7.
KC<a<A(,<J:e7[Q1I_X4^fc-GY7\?;FgcF4O5#O-QAK:WXAQI50J48GBc0()Ae9W
;Q^/Ff&TFX5Xg0UYeW-aZ6>[5WMQQ8CQ@E]F(Y6bRX7&^#g78@>=RfKG?a^=L?[W
b20A+Z@^Z5V0T1F2OGBRWFM#SbEeB2N^dbA<EA?HaPZ0]A>O/7QR/>LW6+:G][)^
QLb?WASDH[B)T9f191?SN<Hd75=W20-V5Z5Z<.\?8gJZ7?Y02S5)_Bg8K-(RGY6-
c>S(e=<=fb]Y[F#:gCEL<9+QBYY::20;OfCa4&HedTV&(e.;=KbPVe3_T]X;K.(8
V&Fa7c?Z4>RD8;[#4b#PPeCTa0081;VH@-fD6dMX\gJONJ/Z\[V[8G3Q2YLe&f)4
UH,dF8R2BRW(H9@(QZM0&XE[3]Te51WIMYSWY];75;3<;N]f6J,(+Z?)&0a&4VJP
,@EgDA2_/eJA^T0UXg+;8)^>#e<T^(5g@d;,d,_YNg.=7_eO2SCc;@O.]@N?#ee[
[(<+JT22gDEYcaV,_1C?A_T(+[65fB/F;b3=c7Yg#RE/+)/LYD,0(4f+V+&e(K9W
8;KJ=AFP.3O5^SceCKLA-fVARP#aQdEFI:HC?W@,1U>-P.,2T]7f9IUJ90I:C7,4
=ccGKWGKR+ZZJ4.aUc.0N/HGP2fO=UQHWR@a=+T7^>6_PI/M;X7ADBJ\MW2c&WUO
-0N:_56AWJaEYaA41&SCA(9+ISd?DcBUgFGS&9a0+^G4A2gZOWf1VB7AKS6XXLQ0
gaa#RB7_-?,S74HWNYBT;Z4<f[;Kc+SXM.K\bbU)9[==6VBIKGb)&05S/VHR]&,<
[,P?=)5WEd.JUJ.\^P=HTVYOB-9L14cP#&_ac_;6LW<-cgQG[JOUH3N;Pc?4ZRdH
0011E\H7(c;Y2[;MZ1RJd_f@33HOKQ?Z4W3fWF6d_8UeW04P.\GKd?4YBRdZYQNg
<6)4B>gJT?)4.5U52@<<R-PF(=8W][7)I-468TT=]?97D\O_^P;#L<MdN-HJKL?G
&TBdSfK?N(U;c]Md)J4NP<Y]IR&]d#N,?I0V02:-U4#f25I=+S4d^YSU+Ke4Q:3<
1:5KNGJ?a@QORaI/HQ[>JR/SY\aF9?W+^,1<DFY]Z9fO?HfUa&C)8.aM31^B]5<J
F\1L?d<,I:)M0HN+5(>H5,<30Fe_EKDb(&T7>ZWMU+LZ<E@E0SSc^VEI0SRN2)RY
7JH/ga[J#4^_GLY1ZA#a[?2K?./e+><^bgRR#J6M_CR=XHKKNa]\IP:90Tg:1Rc#
JM3O.(S]9(OUQ_?/E9SJ54N88f8,:PF-I]]=NL;bFV7U>D.U2bC.6;GL4DDG-;/Q
7S.eHE_Z&9]8c+f4GbU/8T@Y,-HU-X8e.J4dD<-:9f^0LeTO>?d_Fg:P-cAXM6O/
<33R\T[9+dY2@<64&GT6UGZgR6+AU\B@MJVG5e2\]9KC-B,Aad/V1^T_EZbT,RM.
Y(U[eV<:4/]#gHT:GVX@:^.<4<FAFAE-(\,H62I78WXMb?b8ON[G5+;O@K]30A+[
EK+58=d1Z=S/?PS[MT\aaX5,b^QGS;JZ)PMKFd/LeK-IcL9X]^;-\EKQJeO(#5W.
D&-VQLaU6+V\WDZGG#,f-Id@8KEKEL07TdN/\U_K->KLP3Pc+3LJD(e6Md][Ld_/
eX8WY+_7bb<#&Z?SX-A/Z#Q0@g\=7&f,8cV<)L<5O;DAUA]&V_WCJ=ea-34>V6,2
DCAd,VPW]LaG52@E_.G6E]bCb;8-]eCQ1deJED\UZZ60U@BCa3I#&&/6cU&L,.BG
KY.EP:&F,CE;Y]>=g7OI26fWJEDAERUUDFWV&/X_MWHT0(1dYB-7Q)Hb8]:T#[K,
6H5La/Z/55cae^#,J8aUVfT?cJBPRb.#/#BO4PXOOWI,KfZ7<bQ/-/^CGY1:TXg7
@/OIc1\3N:I@CN<1+&-C;?Y84=^3?)38J-0PCDeNE?-IS)V_H,36;JRB\)b;Z-J0
RL.N;^K-F>U3KICZ2(9[;+8OQW3Kf8IZ=J&e40.\89Q=0(\3:&eS@O]2S@FN2a:R
HcaEb\=W-ZIF2O6]R:R[JX@0>W41J&+N6,3LGBgE:U0JWX2?M4Q32NJZfXLI^4#b
:Z>BVWMgM:ANL-;D:)]>4)fZ_SfL.[AM6cb[FM0N\?&(cZ<WFLL]ALR?5]EBJ2Nd
89-K>bSLTI#ddQZ38f_+54X>IbCMG2\e<5NeAXUWH.45b4<?L+.(,E:#Ce6B8(.5
F=U\MC+e^3e_-\VS_:Y/Nf:NS_0dGJ53@BZ>^a<Q,J^?R)R+PXCb[C6g>N\SY:2A
^R]^#6=:/,aXPFd).E(QLF[d[c?Z^].1R1=P68VPQ.++PFA=)Q.#DK-5R?#Q^K(T
COS5C]8U\)L5d(;J]gZ+cSR:0KTQM3@PJ]I)4K7W+ZBdXK:1f52g#8ZXLJ1.Z<VG
I#Ug2g3JYZ4@ABF&Z.EAdKAZ9cK<JD/#1I3]FUV,bRA=:2PJ;5#a2\\72@.3Ng1E
<181_Ib.gFUdS4Z?8#-]c7:D^3UD&eVDYCe5;_\.#W#Xf(B]YQDLeg]0-HJ1G&.0
[4a]V<5]+91C,;WKP0TKJ-d/\)W]4]geVY1:T/9.,>>]cOAQfE(MMd[DVXU3OHe[
f:eKA>N=_b>Y4WRASZU7.c-HCV2X,WN_eUcPO17>26JV(.XNNK(9T)^L\[#<>73O
\5aa(SR+[?6DHTBG:TZa.N26XJ8Ff1g4(<ZGM]\+=IUF8]3f@WOVcL+/8_F_Cf5K
U\J\VH;0\,S-XG2CT6BLI4_8dY<?Y+8ZYDGHD)WaJN@X@XURU=2ZR(9^Z.::=[CG
G4]a^)ISSLEN<_B][)C[A7M:2@855B\]U3\6D/?/&[aZ=>)+328&;1+4DF(]?AVO
+?FGR(Ga1_=+[S;7NZ=\?-HdA#XSE2Kbf=3G:],U9HTZIYDbf<>@NM&[8Q9I&?]3
3b_M+/>@Q^R=a[>5])6>W\LS2f&L</8b.Ob>3/bF/Ke0)6D25^b6b28Bg2V7XX&2
M941AWfUQ^A+-P;=A3/,@Wb<A5J.?YO)#>LXT=EY61@bHPDBKaF3_;3+:M)PFb#=
:@=#@,Occ\gC0SA]0H<WYTBM789N8gT]R&d2IQ0;]6-gcCZC6_,H>N(6,UcF9SN4
ZX^+/NSGD@7)5IS7g6K3VB7#5P&>)7RbE(I(Y?):P6:(=bZ8+6[:B9AO@;_cGU<a
bdIEG6#Q-d\Y)4[JI[P+KFIC&-(8;@5Oa(I)@FN?[L..=MW8)faKMceZVUGgCAE>
<d1??7eZLR,1Bbb2)HP#/R8?>_C95X]b70(LJabRP>:Y)F#FX^8O_7=BFIX6G#)2
UREMc@#QKbG&F8/_eKK9<8e>9\UKY9Wc(egB9CU.T.g&T\:=@g&cJFSdI[VefVBT
:5dOZ\JJa-3ZU0Y>8),aE]=/EK&&Ce2&&X)[,3OI[^O60DV/E[?2?RHabI9.Y1XW
QGD9ZR77TEH-ZZ=0fVMQ_LQ9##PTd3(FFCMXOK_bJ4a;<a_1=&;C+E:OD(C;^TRY
(Y-;Pg<>C>eL7SK?AW_#:T\R\0,\@gB+,d[/>U/4LQa/Q:a4SE3,]a8/?7.dBQYG
bDR^5T9@;J=/?cTN.;&9cdd?S7aKg_.)TV)J5/G)fT++Y=9K\Wa+8&B:N(<QLUZ6
7@_CL57JI#V_QFSd44)=(T5fOZ[_8F9H0KC8OUOY)ZdF]/d+OZ0:(J\7Z@Rg^Ne1
V(X?&b8?]e1F0+JT_2,FRgI_]d:N7eQ-?U1Sg#9V4L1/=JU:_7Y_6IQa=_TYWHL<
&GSB.I=-^:@a)9C58^UVMC^F@D3g\b&fMTNO^aT)E8C]A7BY&e50dQ<AbdL-5&7b
ZYMaL(P<Ob[dJ?&A&Q=6Fb+O6[#7J5U1cQ:P+-)aV^#81FQNgg><L_KcT&OSJKG0
1FO\X)PK)MGbH:ASR\4[18_>YG7UE^P[MBDf1)S01\F7:fKTgF6UZ5W41cYc63S(
,&Z0S(:U2CE3X:2]acI_(ReddG_-Lf6W&>M;CQb(YSCV?.W+AW2OC&4+>H+g:O.+
R>L;@<U\g(>(DA_EDOEQfO_bI9:0E.F/LZDfAZKC(Ib\/N\.2]QbSPF<^geYS7I+
JFCSe^]6,?R;9\[^We&J_&P818gKH1]2\[M73N(cdJ(/N;M2,DcRSLVI)8MAgUCH
T_KL7f?3.g8/46@U20DG_68],GF7C=F9]2]CIE;(]UC1O:5agRXa=+-?/T]bO>_9
bNNW1+Q]W@7-dYG71a0fYXWXO:7=^:TVd37a=QM\FE\]7faJ+?N-7//5aX6B3>@A
)E,NBc7T/\]WW:AO.fUQBR5,.X9d-?QIHZPG4[EeI,,165E3&N5dXc>AY[:S@2V/
Q\e\&B/-e]I3TL#TRB:MPeY.5/H]XU^62F046\P3@_XZ>T<dJI5S,&e6UgB7GGP6
UARD;L?NM>YL[2[cD2]BAbM5VX5QKL5XUbOURKD<d2-[@KRHL_G\T<6fS:O0<4)O
f71eOB2A@ENDC@cZDEQW1;:VKW4[G8_1=>^g0GgISKZ.TTJcbGVc.ZLe<BcKX#\6
=dN/)I=W-TX3.BZ-M6Y_KKNQ6Ff;ML9ZC.dCCCP[_R6BL)PVCYXOf:->(3RBGZ\R
fg:<7HN6/a\(TD\I(8&ER2NYa<1,6<b:gB7OJF;)dWb4S^DM_6U:)+\+XgIb<8ME
L4Nc1.8SROBKXQHX(_S^BI)STa?2E6C9W<LaK,^g4DK/8:YUB?feFbMY+FXde,\c
31T#EZ-9b[WC0YUD0K^E[H_G3;14O]g4P7FW/f:UQKSL.[IE8\7E\[PMN=f5N?[:
5B[c8:,=1RcB+JP3.XGeMI4?W+QD0<Q?Y7.dOXMd+?1/f^;c;=XVNT@?aVUG2H;#
SD<G8&d5/E)];/)gg_:W(.UOH@6cJ;U\>,E_IOS>H^Z,F@8#bG08f,(cTJ+/fN=Q
TP?HW:VQZ2<U[5];?>=4&AB>@?;+=1\-&>:=cHU=&018K5Z+2_0\<b7#GK<I]J-D
5D920\@&_?.Q_:=S+)#bf=S8R9Db3?La<79UG\,.4,8+4WR4VRJFY2OE6^S0M_=4
8^d(XF:1KJA_</7H;\]G[8CV<#[RGDW2RC:1+f?7@WV^XQX#@17C(;Z;dK,+.H7:
[^;8XK#-R]+O=&:-Y-RT=+g(T/[Db?5F+gIWc3S7:8TPT3MZT5.0-7PD7\7-8NXQ
64a#@HgRS&GPXU@f7eX<aEH;<Z3-d@dSd=a=H9e/]-X=+DbU=ISU&J_6_e]AYW.)
f7B^&:>&IG.O]cJC9L[X(]aE=,7F@>QG)QV1gf]>FG?>EPg\f?V_e\=3gBcN^eF&
H3R&)WUEX)(+7NPf-Eb=::TC,<C:U(C.e/Jc)cP(A&/N=DP5IZ2eP,Qa#;9/+TH:
KOV))^FG?,IODW;DK,/CfO]MN2FM=/W/>Ga8R);+ZWDdN#P<?/SNg:fS;(7+0(D(
1I(]:RV)d9B.:N#WOa03\\M)JCW;:@J]dKf_:6IYcc?^5(:X_46<;O/Fe]^6FWgL
T,TX@^AKgJS[fC&:LV0abNJgM:F\4eK9<9_cM4F1P3S9f^H5ZE,:WeDZgHB)9#d,
K+V2_#M\XCZ+AU3,>Q/@4-KP[0EH70WB&BW.@9#J90eX]YA>3KgG[@34#_//(797
8b.50@KG<G8C?+e/Re>?N(:PgP<ZRL7M-O,@V0TD4+b[RLGE(.@8TWd-WLBQd_6W
8I\@<P7-_US+BLJ(D+9BeDK0SbKaXEQbN&fQ=L:LeLT)A9XcK\9:PBIaeI.#gTE1
9RARHL=L&N^MfbD<GN_5EgOb?[BgNHJ3;bT.@CQJN,FI0gX+KRgE^#P8^^fVCK\A
4DQb>R)g<K&(AKSZ2/CCbdFb?LO+PT.gY:58e[HHX)Ha[N]LRO<4IY@S.\<cYLAg
/X&fgUGMOLDEg]U3^F;6YaeOT>GUbf8+G0#]Z_9a-e[_Rf66:^0aP.BgD=0U&L@?
Q1<G[78/N^5[;#N<;.DL,\3fd@\SJI/-b/&c3e1L#HOWdZ;\e\_][#JJ[\8[9G+.
ae,S(GTR.d18)&aFUcU4VOU9QVZbV.Q0H5_?THIM]331VFGQT:3Ra&b.4J\JC4I;
,BRFT#@2QT2^7SJJ;^f/)PS/FXAIB(JaWSP)8YKaV26)KdGMUER2UK4JQ)ZOX,/0
1^.EA4FL\CD/K66=bRcY#@?,-6T@T.=-:_\f+H(^U:#L#+A&g9Z9/S#Kd_dUc=M5
19)991(.2P^#OG))HVde:]C:&(a;f26ZD:LVa0,BFNZ#,bGQY1afa:L[CHJc&\-d
_M3Y-PeAf<UNJ8]W(#d.P6-+fQ-)1JFK8W&-W(N6JR\]=#b/3(fd\LfV^,-^;E<P
?J]WKW]<<[S.AR(-:Q)SK\UY7ef->O=<5BL/&MT/5AN9.+)P8Q&C;C1Q>25PVUY)
CIG@Tc.5[A0G^C.GHE=CP[AF\0+-5535K.K8#7=5J(,&#e>f)Z:&PMH@F4a9a0FU
FdKZAN=#3;N?7X&1D4M(bM^]6Y5\a^#\a&EUCJ;BYE^\6-3@7O,J/GWQ+Y#/Z0FV
I141[;P5RdL9<YR)Z=Y?Z0<cBOC-9QT+eX2IWJcC_S]M=1>>VdEbZd]#Aa,FMIX)
DMG,?+)USaI5_>-U\60deO+da#Q<#AS]CYSM/dCcO2IJ31MGY,a\PZc)f;Z1e6&9
_UV-eC=DC35Y:J+J[_1Cgf:]N,Of1<#AM=5T5Yc=#)3F\,He/ZF^eI+Z#,O2V8Bc
RAOZJMf7Fa_@MB4)((a+b55#H_G02TLJ_\-de1_G].YTOQW.ebXd:Y.Y#M-2IWP5
cVO&TFJJXJKJe1SCRR@:5<XfR-W\>N_<GBE(\-=::&0^e9QG&&e=>A)9/41;@NPc
RU2,/Q>BMRP=fU_3W:/P&G?b(F;P-?<DZ:?,g[6>C\N(O;))W:-RTf9HRGO(O&a_
4D3]]E.<:<?]aIeR3N[M\QS_R#).QQDC?:<2b9cP_CDXK?a=dHVa(&UbDX9RC/IW
-Ud)eEI:c;?f&(^Z76H5800MB3:?U_fcW,T6_eaYWZ;CefZ<A0?Eb<>&a)]XHd[G
C>/AYcXeSJc1=3JX^HB:AHdWW#7KX3B<8IM<EM1T(9>9SR2GEHg)(>f-4U<2Z<\/
EUd-GV/=)M\T\L__b;g&3<@.Z>]QAScd<O4J?<W),.dCV6Tg9(gIP[3?#LO+653e
@T?VV,SGK:I,0P#].ALA-(_P;CY+^0LLC&4K,dERP3N]KESe@,CZX?3.AfBTEEQc
c+9,6TaEPLe/W54\1.F9)#BgF:/7ZW];XVb;ZI14H9EZd96T+U(;Hbfb#.aW\g;^
gI#V>((G;[)P@P\T-gDC=,KTK^4.M5[2)P9>,>-;J^K?<N.G<=J0EG\C=?K:_PA)
\JX88\6IN7Fe0F,Je_Y=@T1W:WB@d,U8FIKW-M9\-B<4V1;bcTAWIOfB1-XK=2[G
f,1:=b3#929C;@Le.]W9F5L7NAD#H:Cb^6NITA2GePD&B&9WFAE@LdHg[#EECIY0
#MN8IPC/&S,QJG5LY[DGYaKce/Qe]Z1Xc04gO-)g(>]YHN7cXc,0dD2VD1]\SL/=
R)?ZU_YRM,/Z,0Z:-[)^gDc6dAW]F^,7bc0#+JW(15,f3L3B,AZ712eE8:5FDX@S
G804:<\JbH[.1U8W:Q[gdbA\9V3W-]HM&<_/)KF(F_H,U;:IE6.TAYc],M9=L#EN
NIaX>;,0&L0IJfY]>R.R?R28;?>7@)6QebJK##+^&;@>-HSE(8RV+=>U0f)OWa]A
=1;a1-48YD5-A;81>gKI56:T23f,S,/_2VQ]@Z?SHF?UN@A&X?KJ3S/a3#JB]TN9
3+gZd1DTR5)Yd54(Q&]C@Gc>4C4L88:dW4(b5dCHO)17DSPFfNOV:O9EfcR,[6P=
;?^aH3-V])F4+U#aX7Q#=@ggRWW,^bWcc1A7GW6/AT[cL21--PDY0Sae<bNE25:d
SOK91LS.Ib^_[FeNaRQPSD8QL&<=JeE>&PT)GFEg+9JI<07)F]UIdVQ[+?)baOOd
>V^f6^+51[>FR[AIQ=(C+NAC(@L=1R_5][5=K&1IBXIIW_E.=LO[0KgV9=&4@9Y3
?aR27A/-6;1_5bX:N@XEZ<R//R)SdW_;<d[->dN@@AY4OD#:F?81H#]P.YWK3X)3
B=f7:RcF<9:M@971CcfbRGQgN-e-J>.LT1<2YOaW5@]1H7Vb9M:CcKAUQb+N4g>[
Fbe+Ng^La7L15]\gg[(SbJa=ZeA,F<)+XT5\9M4\cG(:89PR^9W^LZXNB++NP6c1
O&-+Oa3cY-7)00R:)7L]R&f8FDTKKg^PR[+3D<_G=^MaX>5^]K472;H[3#=?/E-^
-4]Q_-bPJ^Sg^F40GNG(EfXEgVc+;a9]dL7&Ca5f#8+&:5CFJ9cC2O;:<)AWXZIa
T,c^AX(<])W94C,:JAF][/G3,H/S>\)&]H\@GCIPN)@F.;;bJMZacVKBB>8ca:3.
b+V0X51\P0_HgJX>@@,c.E-B4216A>ccJ+YW&WXUG02ZC3X3DL-ZVWgd>88K>8Nf
c8=3NKdPV;d\[bCg4/5\=5_[7ZKBDbM[Jb]F?6RTJ5eb@RI:a835MT<G1+6/baRa
;QF]8G\>62KG#4C7?7(#aB)23E>Dg0GBc:80FbUP)1>bWG=c.8faeFJP@Ze#UE?[
#Z1gea[C+a#3PQ1fK<R;L.WJZ=1A0\Re+3JT6>LH3gV[)(d:>\CPdZ@&L/8)X+RL
Q>N>HX@Vb,T++-6gKX:RFE(aDf[BQ394I5,?.FKWV5X:7g/P,_K8#c7PIb:5]D+O
bF)5A_8(c=:Wd)+D[#>5H47Q3#@>FH(^YK>XNUAa/BKK,GN([@//6S.=I-_R5G,-
Y_a(d+F-ACg2_B^FbU?2c;[@0EBFKc:56RbdZO-(KH&FLaJg.@2bRN7[[V)Q&RUL
c,T8<e(E(5bN]+D-gWA&gL)SIICK/(Q.K-cdCKK[MP^b1QAb?0edg,,D,BTCd4C-
b@S#7T94/-:g73CK1Td9D9?+DVEY7eU#Uc#FO>K[>+[-^d&2(R:3F=A=?DT=89MR
A&?aK=I:T,@12&TM+M07VU-gN_Q=/LMIF@@M_P?/BL[ZYBD_J<5D6[:A-95J,dWc
EV#;2+U;TWU(:MZZ+6[b8_g0N3\C7]ZcUG4<J&>\SCEIA4EEIUYY=bKA6R;+7,6/
8FI@6ESeH8+LKB^EZ<BLU\I,eKb0;M2M@0U03c]HE&O68a=<>27AQW\H)SMR_PD0
UfG9@?3\:O;-HCCWc52TF]9A9M>+VUD0\0+SA2<-gO:Q=(aDCN+4MRPD7X]W>G20
=;6.gLNI.^[a5JR1WFA)2VPV-23P/RJY7AaLK8MKU6L^TO;dKTS(U7L\W4GR1(HQ
NP+cX[O_+MGI:?Z?:Ba<R_OcZ/R3fKd2Y#:JMS4LS)UA^0/2I1gJPFXHOB=TA<5J
[LN>5H5bZZJ3B5T^^&J:H^KgCX?UL+&QLB3dGAOVCfU05.&A30B02;KA5Z,=4\<5
^?/d<C?2<FTALU^XJUB8O;P+9AQgO1C5BTVUHeaNC=7/T\\.>CV,62[V]18/XP-,
A>JPEKV.afL=:QR@EI,c<6Z21W/0:)2RS,>ZND=X;U9X0>3b6:0-J\>:LB<Z]cR;
F<dN4ELQaXg>3;/;^4YA@TN32OLcFDH?dT;7NXGDXDC<MdbA1FXX5.:Q]NI^SFJ<
_+#(,R7f]MVY)_7F,/6IYTZ91AQ1.WJD617K=;faf\(+a3<)/HbDP-ZUYdNLcE(S
BABR:O/UZH:]9fU^)fcP\KTP[:&gWD<V9VO,O<XbOa-9L+b^?2[ZM+KQW\\1>.BX
8H#K9?5.K@J0b_86DZ3_H[;>+7D2)SP]LJ5,>VMe-\FATIOUa#;e;&[Z2dNCS3GC
0<CW6Q;MC__[;YA,AOQ>F,EPTEaZ-YdN14#B+A._DT#3dPN)3@F4CT;UD3X^_b7T
af2KZ:PAOdUW#ZYGL9BNE7,dc8CHcSY1]&5)\J=+UY-GNQ:RaYKUVZJ=1+Y6B;()
#0T=JUD&:=TWKSXdB&<,J+b+/c^5J]XJ0)4c@-UT4A8H&Q]cXIB=c4GAW?>:4f=#
_[T>e;1.DF[CCR(W07NF896MM=9DNSEbb0)@\LAP&#^#VR1&7OLQ6FW/J;2KE044
PSFcKT7]dD:LEB5J^H<DK+0/+O7RZ]Y>E1WMBVPa(D]Q5/43JUVHQD<^P]L3/4QE
J;-Ga5?<OJ\\_IMJJ5[3(eddO;?7S^6/;XQQ1YCeZ4<aA5_S=>G((9D+KWL5SL#A
:DLIaNBT/e-P2I3;0I\\FVN@-.,CC;7-,bX\(6=JKB0<_ZDTPF6<39c^+C=DSV#5
:KeAALL+14\8<5J[If>G8L91]bY)YQA4aCAg3+ABRZcNbd\d[<AR8[NLV74UH8SV
N@0deaS7MO)&D8dT_CSWUYR]SV.D3eeVM-g^=<g:XL=VQ\,CERE.:O\C7;LL4,U5
gcEH3AJE40TYC5Y539DRUSMF-6AgTd2Q\,/@\=RBK6BK\d.#.\K)Y9?)M@YKJ6<H
6<]P?Ka0]@F=eb)N>DGMRXUV3-(UQBGV>cLUYbXG2=P6:A(#4I@b4FHd.9M4f+[F
RB9.0/?0P7J=?Te?5&)d?5L=NMZGJ+[5#+-4,,<EU-LY-Y.TNMLGf)^;BSF:(,VB
>6N,SW0?KSf<9QGd@I7)^cW2g-M>AaUYF;?9X?H,#YF@MH&00\G&&QTK<A3MK##4
Y9b]Td/W.32WOJa&5LgXS?4/VGV-E=\:@f.?BE7MT>LU^<@I]c9BW8@^dbD4+_b<
aA8063?0DN5T4II4SX:;QDcd=gN\):N4KM0a4\=DK^[Fa6EgQJd8RR13HX2O/Z:>
b8<Ke0fBZS-0)G0f(S(S>+cN?YN<65>];0Ra&4/AG;7?^RFE3O6HC(IO)=3HI(O2
TZC<<\&V8,_4(9GfQa5,M]:.O-eTU&6SDQ5.JX\2:@<X)VD[(<gQ=;FPNJ=QNZS7
W1(/B:HFD1Lb7X2K#7f\PRF=TF_7Yb8GW2WY&AcI=(-;,5CUHa24AX)F^BKA/^Qg
6aD/GM5DbA@DK\4&G46\WgA2.39])Q?O;+]gMY6;W2Q>X1?@P^TCH)S#4,XQ>R08
7HYXX3(FC;^5(_53?:Td7fE_bQa&[dI=@ObRC?#[H#5_[Q+#MKP=H]CT<KA8S_^>
U<?D0^5G[9Ub/??g,M^^#2-fY-8F=2aE@8@Z_2E136f&0_+<I??P0:_A[SG3d[fF
f4(&eAN8EbeJD_c?YV7:H(FI61dgT90?RV2JcCLLWXH7GDcMMc<2+W9N&TGgCY[+
cbQR4JKH8;a_9<Z2?CD.P6VA()Y-)JA9e5U&>,WCH]1AGN4XYN+&9+G@CK@=.:DO
OGDY?@E+Zg9O/+S03?HKIXDI/V5R?YeR<O?(ZDPSXSdg0eT?-0)aV(Ma/dXUMGff
AM2D=WAcfT[e8[EBX\A^X5eW:JB,Q?:F/L>-]5<gZa(JVN;bN3eGD1@FEXAK9UJe
2LWFNaT968GE2F8PD2UAL<OP)Og9IQ?^>HK./F<Vg799UHd/6E4MH7OG<X5X=-1&
\RK.;?^:N[NS4#?-I6+AV<&e5/\eUAf1<OdgN6)FYZW37Y4dX5bZ\D.VN/U-&gJU
M?)7F]G4Y3#D;_[8UCYdc9V9R?.WEG?R(d?3//[c^+7G8(HJU<U@[HR.PD6A,7-;
FHdfQJ7Y;KGV6cZ9UZH51W@+b815.+3+==W5]fc]R463J2BBW^)[]H4Z7SS\aVTU
_Q7A[(5X#.e2#U<Q<Gd5e#g]9O89)e>gII<e5F:KdO-K&H[gQa,6O:DQ?fPbXg+8
f2b(WJPU41OUK,UA]3]Q,L8eN>1Q@H4DW;D3AVTF8E7fU.3,7:_PV=&NHUb1aQLP
&=@TZ\=VX-EY-ISPa23#IJaPEELFDbb^O@])IR\Eb6/1gO[gf[^OIW1I=K(C\./.
[7Be;#^X<(]9#MPI),M758UPW(CfO21egP-HS8HRE8,4<SUL?DBI_Y),I4K_;bHF
1/.VUb#F5UG9[X)TaJZ7c_1T\RA^cZ/HMR1Z2KgT?e8,(J?]F-35EB.FCOW7FC>@
^3+gS1O9=(G1])[:VAcNW9cI?#(ICKTATG,<Pf;dH:F9_^/Ra7OVNg\?:[=-2R@Q
[cYc_<PK.d0Z,E>X[@ddYI0V<Y+Rc)E,.E<Z+-RSS^BgdW[L1H+X3L1g8f3+a7P3
73C2W+^dAP@4_W5be3C<?(HA3K_7V9,(9Q1O<+V;CA4^XM?@8Q8Z6[R^b\XW1U?N
EVIS;SNB)4EXS&<CC^;8]b<32O?1&I>/??=P2-U;A)RP:J7GJRR^c7_IV^B1Vf+B
>:b2O(4.ZYL[M)bFHdLI=#7:..H=VbA5([I?J0KXEQN86WGT&JeREXU[FR:O1Q8I
=#D9f.:JE++:DRR^A.5X.+(D_:E3<N5_4UdXDRN44U9MJ:HaCTNYHe.EHH5Ig6IL
ZLPMfH(He=G;(1W0_eS@GQdGc&T3I5JYPPA:I)\P3c.-\(Y.gF(E>UA7J,[K9R37
)1?CLO/:Q-+[XeFPPTOCFZfNK+^<eJX-VXI:Sgg6S3K?,)^/1aE6?,H48&4Z55<>
V[b,/GP+B79Y3,_^d6<+Z0Y,V-O-C3.Na_XO0OV0T7NCda(NU;BgK2N)K7)LFZ1Z
W#OaU-e0,9NU38CEM[B9JMc0Y0e9E#b#H#=V@66R5Ec9N&J<[F4_UF8GeT=OU,+N
Ub3c/]KZMC^9IPF,e(](SA;_^d3X_??H]e+P8I:.+Sc[BSU(KN.)C<O3+HFG#,TN
c.Y^&JOJb^KddZH\P5Rc3L_U;]AIY&(E)QTBL14-\ebUWGHKI[WK-G_HA^^RA-+X
+O24;@4M]PL8YZ(;+9/46gG\ebRV=C@Z0V?f.I#R^;Z&&@;U#4AR(<E5)XG>;K<7
B0DLDA46,/G,^20&P/X)LQU73CL(UJ.VVQ&c@4a)@7VW-/\7V?Z=MM3-#N:RBL;C
PHJ[,XG81P.[RM?M4D<8Qfa:?[3NA3^LM)+F-QMa<PcK&VB7^F]2NI)L]GLRM=e6
^AH+)#c,#\4+7Lg5=X4f+]2(+9Xb;LJ8-BCVa1b?WW,5+-#(b?0UTdQ^fZ7>/0S6
0^KDQ(N8YVD2c-@:J+X7:&fYQJcf?_)e<>E\Re#IdX?KA[53aOAX>XASZ;HdFCEV
#]7?(3]&CfSWB.@0RTaPdBF++H?Fe]X\@-MX148.@Q2?W3U&;[I@)a69AQ;L,F/A
3O@R#W^964[>I@C>J>/bA8:)UDG)T9C<TJ\__&eDJB?)+Ob@@&1J5O^D7IKX2<8D
N(7PfU4cD7:.VTg?CF6fM&.c<N47\Z]^<#=6Q#8LYPc<B&PL_(Q5H]1dME<ERMQ(
Q+c>>OI.]YG(.C#D#>I:H+9.?<Hd5WI_B]ETBAeb6T>_aVfe54.[7@L<>,2;FJ[J
TaC7?#-Y=N-He>C?#^_64XT@VK#?8,E4N.HO@UeKQ3,OV=d/a^>3GQ7=9;U^&#Vb
)H>Qa@[@PXB,bePV.[c(2L2-,30K?)E&eZdF4++\?DGD5UdSX0O(F9V&2T26MK/#
X;@gP^[0O3JX?J+3?]14T^^1HSYT6,>19#];9\@CceOA&Q8eUa6O[03U&[LWA#1/
Pf[HOE(5L]+=b^g76G_)8#J#I8ABAWEU3_c\K8<[A-=YC=R>d.OM:??-G0&.HC5A
GW9<-TTV)2-PE:63KWXQ]WV]&T-O7fd.?PCKDJ:I\d[5HY#E^CEC)L2G(?dadHB1
G;<TZUgDVD6.7L9Q6:,U_>]:+@7/A>22ID\OeDRY6;a]:B\0/38-W]P0Sa?;Q3V_
B)5N]CdX.YB)F2bH](O&GU&H?_JRf#DD;I^4RfRJ#?&WOX-^b/b_g9GT:DbdC98\
(P8gSA^b:cR8H]H7N5/H+Q74WaE(80P3FA/LB5GAPEL7A3Zb+DN2?]>.;5NL<ZQN
@6bBZ,]9FaS_F5Z3XT+b3[C/ZbG3Td&]Wc4YcLQ.MF)R/GEH_@QF)K6TJ:>P1XQW
FRHDZ6XS4+](<LeW)<7E]E0;Zg3EZW1^5W+e,IM7]aS8N5-02&?YbVJJSQ_]P>;g
<PD=-&Zg]&);2S3HL@V9?e=[YZ<?5S7AP6g:44S/(]af4)@OdX)Lb/:,f,[[.Z<D
^70=S8866/[WSZQ9LXTX]1)FG(58ISabN(0U6W.)MTE4:ER@,c#7;Q&2]Ka<1e:6
2K\]=K,;PFE86aF-XO-^;MCJ8;EP.;:3MM)g0f]F39?<QW-N;YPg4:CFI-6P:RV@
@L_1@(_DRI.PB2Lb?GG?P3^5K1\]eAE_BUY@6R8)S\_H_+BK=53M38((+M\?4fD#
DGI5a#Scb#NeV9(F<9^)fG,_1:#2/^L:N&L(U,@5I?.A>5gP3_N^[C4P1>b+=BX2
PMLY&,DcNV+O\@T.6AXD?,[C?fB0SaET-_dJ:K/bHQa@R06J36)X@I=P[Xd.E+0C
[;eCQ>eXACdTI023Z#e,<6DBO:4N3LT(XeRB;#Y8>g:c;VWb#37=GaB3E-E@TVMc
;Qc>Ac6H,QEFHIW?)2gRA4M[0PI+-T#MK+WU<eBH[6==Q+f]=\f@Ka+US@29+6Fe
MM\D1]@<[Y;3bW6T9fM[J^#X)7];Q5A(aZ5V1,4ZdH<^YC>7LA9YZa^UR\2/L(TJ
\.BcTEX]/eLK3AEgW>W\MBcZUJ8]eL&Ogc1J?^D4ML2LW1:&((.47L]01>&SB-/P
HV1^Q(<YBA@-\V,&3>g295HB#(]A/FX(HJ.29<MM7B)41gVKH2bbCeN\RI3f1VJ>
-Z3)BZZ2a:41QM7?^Z.L^dcB9]&g(X>Q#EceDeXf@f[X#FELX^]NeT5C=JC4H#Sd
2RT?O#2F6BHVS7NO>(&=O24@);PU?.<O3E2;AH(^F;]NZbQ(=K=c1Y8CP&+CD.:1
E7I\<GSL8P0&IPAIX:c>YbQ<Z?:a40>X<_f[15.(;RGO>EV?3bb.I2@_V>?+Ag5g
O&@.3/(Y6F__H:S4T@@7;8(;KNWf0O20<W;^ba)2008f<>#Gc[,[cNAFbA>#b1FC
GY?dB,[T@]3UA\0[\UIM#\,^aX#e?XDbRBPO1J8e3BZbEYN)N+V=ba/Y6GVb4JD6
0gIVS7)LEFFJ6LXfHB><N9ZeV2Ie<@;4g\Z^HHQX0Wa_Z_UL9@L[a8JVE^W(Ge4^
:?<IUgRAERU;dO(M/>PEJY\=ZOWD\7&9c+3+YEUQ0b:Z;4A18;&GcSRcE07YQ3O:
A?FYZH/:@DVU]Ig?\@a1HTNG\XVa@:<c@+437>74I9PgfW,a0a6)C]bf.a)E6eR-
a,,?6L#,X[A27O+LN\8_+fSGKD?RB])Qd@[X+^G:W(=?,UB)<)BQ;M=LA3WZL?JF
#L8/S1NZ0.M_X&H[H20HeUZ7ZQcZT/&.<E&P&#P@Ia]-9(T/]EV,gB^Tf?(bLVO)
W)<&]W4X9BNYcT;LJ7,GC=JMZ+Z72g<]=dB]B02/MU^)OHgbBHD)bQ6Q-#8-#Qa7
,&Cd.4e7D<X8Q+3dI(]V/cfO(PK,U0S>Wg,E=M9SMCg8?EG)f=ZQfP5I96:C.Nc&
].9KNc-:=)J[cXRK&DFA>N.9ICEe8/L0bYT(GDDOA(?5+=B=R<@2fRJPMMRG;O/1
#??e_;[-XfcaaX8>3?a/(bc38Kd/E5_@dVNIHK?T<b8\3C>GOba3Wg5UI)CE&-Q=
@-;2]FKHA\Pec(=D-(BG^#ME3:>UN4XP,eGZF/:Z9TF4..?Oc0_:88^/\agK@P2d
Sfaa]UQGI=++/Q8^FTXBLXE8D@FWQ1)QaO>_A>cb:AKc6@-UEeC;]gDJHMO_AK1L
&2&^3U+:5@A&:P7LQVF_(,V8QHH??P=1A;)P:_H\C6dT8\XNT2+IW_/@5b>TT_&)
G_[]UJa>NN-]QA#3C9RV0>G6bJF0A8HIP-+=3eLIfDb&bN4=O&AK&eL4C6&M3].P
?[d,.UI0&4Fd0(Ef-ddKQ5@<]fK3#XP=Y7GOE/gMC9c@&#U4&>8>aV?ELd+:#A51
e5@MFP2B&AV3d-_Re9>9>;3dCB\N3e-/-3AKQ+]GFa6M]8JU]Y\K#c;RR\6E6^9/
DeKMNP;fa&7_T9YabJB..aY.7P3-#_-F7cgMC9MMBTgULR:S:KEPNX@[3:+XE,)+
90]U0O5HXf<WPNZ_G&RL_RC)Y;7MG3^.4+d&R;EUX?[B>#99[FAR@.BSgXOZ(Y=7
0MHOQ-c5g[<LEP+<GRc6(<PVXIF7HM-D0[dFF/?Re:5#Re(GPBTZcCSaZaVU&RQZ
:-FG@6T2&\d]g[7Ua\NIHe;K?P3#Gb[bdV@E2+K.ZDLFd&^LYRC_<H#A3LZ14dbd
<fCUAWJ\PbXB#^GOUe0<WbUZT9g+<ACD-DSWQYA?S(/;W:&E6d]g<VDgg[<>RK-#
\QE9:T)2WLYSK10C]ZP^@Z2f&?))ZBD)K=\KZCgd9^3U;1P-;)SYRRbDWS(C&.,;
EV.G92]C0RB0NdFKa#ZU5AC]2\P]C2c2(P18PL\5,&6)UUf^_1SAZW.:1ZE1W3AE
SMSS+LY0-WfA:e(RU_?\=8&7L1O]YVZRMa;(;8/M[AY88GM=41McXXF2K;)Z8?W-
+=Z94dA];J9H@=Y=9Y]aD99O5D6ZVIc@/)VYb/Ta\Y;,6GPTX:LIP@g:>a_c5/#H
2dJ98J9ZQe#=P8Vd0B)LO@Ze]@V7c\d&c0#8BaKA86)g.:N\]QL#@V29Vg;6Se1M
bP/GdLK9NL#3dd+bZHc6A4(=c=-,[>Z_S;,dcNCA6HDP/\gSC?b29<EI/g&6)+<-
RLQ_S7).;CRLI7eEJL3YL@X>2,YG)X9Z.&XU,P19@(W(.V9:<T^Od8WE^)S#9WG_
SP<S^M.gJ/L8PMC9;caV_HgaB/Z98>3KY]b-I6f_Y:#g3X;d=MZ&]E]U4fGeJ91M
H18EV,[_\;Ig]SAI[2TUU-F;ND8[&b;2&@<N?C7>L0QQ>P-.KfF6LAN694]E2\)U
LOH?3CJR+Pcf#(516R@aIS8.B2WCM3IeE6\B#H(:<..E[:R4?c#B]S@F>aNLL/d3
:2#I^]+f<+6QBP5HbCHV&6I)]+(1Ba+>c;YfaPZ^Cf_AAf0_NB2?]af6J#CK4b@1
#G6^X;FeLO_V]a)ZJRFF(K_>F<SQG33SPG<063-^/a8+YJ(Z/cDeWO=QC8PJ,KLb
.Jb8:f0]@-//))D2.W.HUH]C1OD(O3N_YD7F,WNV,:g=JDeI4+O;IbbGQN=U7^UM
9L/+8d1d.SH5QUS+aKK[.Af??#3:eQX^5SEgQB[S,Z769NQD4@PIK[MLf9Q4EHRF
4/V>2I8PX<AF.MSYdP9X/V_dMI:CdfJ_4H<\C;YF=PW9\3Y98cD(B16(HW_LeT8J
DGY@GgI]-D2dH]J[AMWGZ>.4BBRT9,>M<B7]bd^B2V2_-QgcQTgKQ_)[BXEIX@U1
ET<f8.g9&M-8OK_#OKJSE2=bN/W;2_McdVD4]JKR<VMO)3aI3^\(CY2GVHKS?P?e
X^&0(\D68/S83&#^ZF8N73XBRC>V./C6AA\[,.?8]9BGF+g1K)a9YJ#LH(/c4dHQ
S>P7f,W;EZWDK>.fcXZ&b(KeW+_0b7UNA7R#5<.<,UYReEN3e<JSPX+fC2I==9B^
J/U].F@aJfJ=NE9G@;L#Q]N]1_H^ME=/A_X4Rg<c(D1#131-ZdfA:@J3,RC,^T1B
TRA8DR6Ee_c7]b5E/8)?GC(V1S0H=Q/dZN;Q.,&U7(@R\W]fd^5fZ40U00[[;LbL
?[.<]/33bGBKg;Id>R[G\LPc=eOZDG@\Ga_;Gb])N1_RY;4dU=M3cTC7U)19Vc@L
^W7NHc3.e74e\@b=V#]\e,\;<O1FT/.fVZ@6JfC>>A3D/U4^CD2A\1ObOR:=9W5O
:R2XL,8a+Z(I8:B_0=D=8F2#8C\ILA/_5<]ORdV5O>@eC,2fE-VX,N71^2)1L;P3
L+IMV/YH:0;/\F>6Ugf6>Vd6ZWSHYaLVDFQMcXBa@]J;TM,57EV7eG(33a1Ja@M/
6eBeC0]Ba)T]&B;CZG?<M0@Kb;L:.ZA4V]7U(TP0FOZZ+V#M<cbbQZ&bQQSUTC:M
R6W.89GZLIC@,fPH,adXDUX-?Qe6bF0F(48ObPJN[==9-3EIcS,QL(FUW&WFQ:Wg
:e:@3CLZB-3A35Z9KKTS65#\gDJ-cdg]KAQ5W9?GTaaI7KWIL@be(@>6F@[YZ64C
T6]G@71@U1VEQO;XSNa\LgNcf@JX&=A+RRZ&;)MXIH;EGP@82G2#f,B:d)S.ca8L
#(]?00Q8IMf^:.\-E1N7GJ35QB[L6g4L0eT@b9RWV=5AV/O4HPGCYFY107Bc:\7B
P&KU\36@Pd]-5\1U(G9Pc6NXNe3CRKH1J995R@e6K=Z-P=H/a2f&R>,6W8L<RGGM
9U(\96>_BR.[#2[]B<F7aUbVRVC=Z92+&B#60/3<[^UR_.AL905W?O4J@dC#VL10
aJA=#Z[F37g9L377&<^/<JeZ+&F)d?J\A:/_:WPeT3#8]A/f0,1N9bg]3\[FSA.Q
;bY05Q[=AAT4]M;Y(2=T1@-OLMPVXR:b-Ja0cP9[I^;bOb?R@7[JB81Z=MOK7<#g
9\&8YM5S7ePS^f:9Q5T_9]C?,=dF]W0Sg^WV&S]GVfL-c&0N[.LGHK9CN_((B=5\
J0F&2/7Q/aIRaR/4FA&\dGPZ)8+051#^IZPGUILK3?R\3S3Z7aG)WOQD=@,B9dLB
SMUgZA[G?3/CSXT+)e3(ee^G(;/d<J@X.J5+5C4;#X6G^11:4VWL79^]6.MFC4ba
R.IOU^C/@0#b[#5C+bCA:_RHLP-.g-B<0TL5b@KWA8^NEWL^U],M[R)H&1#];WVW
US_2&\[+RHNA?GNF/aI03H2fA^ALF]d?+=S3WZJ1?UZF;Y0#JF.QQFRN:.8\Q[@b
]XZK1?2P4[NRge:VRB3.F(5(<<3W5S8P1]NGYYZ8_KHO06D>-,MT1&]>6d,CMJ)V
HcUSAFcE2W848GG#O/UNUJcN<A_aPVBUX8SYZ,H2O5GDgZEfa1db-#3LB<d8.If_
)NZKTX:]#DK:5I&#T>QH)]6\C7#W?C:N-J\EB<QYQ66DA725NF)]?SIWRQ(./_<H
F_;C4=8RTf,M5K-UZ<FV1=1UbS1LfM>dOVV:]<DS2SO6Rg:XLA^B(D;[-JDNB\XN
YX4DKYV_Jb@BcUAcF2GL#1\I98PASF8-4GLVT=[TM>WHWTGCTEL0/-?:T@GOAJf]
I>A@D^&S,IJ@)7LKQHaZdZ&2MEGO_C(2dV0Le)YG1eAV52LYB7#c9KF#GK]78B#4
A.<5+PUINf8U)84(0PSOf>c>9USb+(Jdg?F@?0OY[@VY;&ZTGF8L6;M<L2AffFc?
)<-CdH1BT5>J:4?6f9XHa2@)IeJ?<)2e4L<3ZLJb3>W+@#cZ=]Hf0:8CD7T:C6YF
1V1FADAg8J#UQ-f17&cTU#cYfA#X,GBWd.M\6(6OP:HVW@LIMZ/MYNC.DI1c;(aT
-Nc[,9JdR^O^c:\CF6&QC-_adCZIRFJcM\g7BJ@L+5V:81Hegg=,&;,80=#23(.F
A&+J;7Y.U<3ER2Q26)/BJ2JS;ABDQeA;1)__0g/:W?S<PW:PAabVWTBE#DJ-f.+Q
^AAM1\D85SG?\74,(_d@;67J;SQU;4[:NcZD5F:f7\7B1MZKJb14FTA:J+LLRBK8
VQNM2I?F(B64,[?7[e6PIcFP#T=Q_]a7T39<f]S#X6LVQWgX-]:LTagJU@<=D_gG
>ag8c+gXXZABJ,dVR(G,)01Z(gAHa0.>HLTfIa9?8Re5C0H>^SA)@4Y.@G6F]aIW
)^-Me;]3g1B)9b&?Q#)fUY6+Ca;#<;3K4PR^EQ;_I038>DALOcbF:Zg)-RL9ZP34
<_.;RY8VOObLPMQc,VGA13AX@L:,R_/a>?8c8[YWQ7?H_a_D]S?<&MH6Pc3(baJ8
C6;KY,()b=43dR/A;1>#H,YY54+@U45_c84ecY;^Nc[U2+HRdB-T9ef4A?AU5ZC=
F+I=ZAg9F+\=I&;ETQI1ZeRVY]PNR/dH+dG#[H]BB^B4R>QDY]W&\BMGg7(NH2fG
_(8gF>([8+&QWF389(cKCG<S]OA=Q,LZ+;)MQ9gL^=6>\e^)3WEPL<B?@K]C1dOG
bf\PHM0a-HK#9&)H4C,RDU(Gg&10<R2,O[7e2PA.W?:T@Q&3&APZ+=a7J;:H8W5V
:I4+0)&E?\\J8,EG>TA7AX;_VZL6Nb@=Fg>50U-A23I8.ZYE1EN3/)RDCEJ8BaQ6
@,2b&L^CG-Rd4+^N9?0[6O37_USPJ(Z)2U&G/4R_LK&Qe::\C2[E?ADYd4(+R-a^
&3cY.R2La/:Q>a\0#Qc;YUcb,AS-31#R-\fRcQCI&T1F+N=ZGM\15g^SDT.YPWH0
9TO[WJRcSc\7LX4F<N([.:d<SNK,YF2WDNG1HJE7Ze7I_Nc9@_c&5^6MK))6L]4E
>1a;]g[\fBF;T++&1CaA2XMY[f-,6-cIaC6bB0&73O\G6V.<E8LORB4-cS9/FE@7
@[4&>P38+<+1XV==8K#]HPZR&WI,]b<G(=_)ZVT9+DY6_M+3?VFbACTE?6;g?0ZG
D8GG,X3E5X40aV=M5=YVX.Y8<B6N[D1;#g3?d5WT_8^=/@gU?TZ7fD=&c?KR6S>8
-.@dZ]8X-VQW05d?=-dXeV?)_&(DMTW7_aJ&/ZSS<WT)d]6gKB=4Y?aNC]fH-F9g
YdXBVS;5g#D-b&D&9FGaGBM9_aZ_]U/S?)WRK)Ob6-F^\Z(fA_20,:6;@/_MCD&V
?7UCcE2UNU)POX[?d8\M3H2.L,(#/9.7,#\E=\RVFf[_FJdMeKXCF&<26g+.g_:#
F9(D2U-<EJDCaN#6U2XDe/3.5:QFUQ)gKfUUdH9]Z]?KYeOZcZ9g\>@O_b>b<CW8
Ib?e_I-BWgdc]<RE59AA_FB=LK3b?F\W/dV.I:()D>/G@\T^C3(XCf.F:ESe#69,
8bZ7:dH:F<gLQ0).Xf6a.OU@G;d7&#016O),IWaC.SKKf?g,3.R[&:b@AM:;^-0J
/-01be_\4_eAO]e96?^3PX.R8IXYVY3ZP-b0546<GgF8TI5)6F(5<7C]0TLLFUH]
HPG4UPD=bB=^OL-X13FIZ=d(+912?US9&WV:GY.E?6C^D4]KfI<KdUNVC0F#@ZO.
^H129M<N4c,cL@UK;H&HJ-#2Z\X7?S6.D\TPD_c(KAUD?2]QENYaFDVP2f3I7Z.E
BBQ7bScDI;YKTZ9\VeA,Y?-O?/d0Tb]EBeT9WcbACQUDSP>f=J^MN8+WFCP,b^T=
ZaQTM5>VQ:6>)GKNRSYINbe3(_QS>1:39MfP7SJ2@UT:H^E9g^d\9-d#Y1=gY7I?
IIQ3bIdFR[/f)5fZP<^,WJ/6A,3EVg8.:L\/J?O1?1HWWJ7-V4@^O.T9VZKa_J=K
XLDCO>cSVZU=bH=32d70L_CaO0]=V)MZ1M[D,PRRF0g=&bB5=TV=0WH50T#5K2Ab
?d;XUBIN[T[<<+[.3<ABbBK);gU^b@QTL#OZ(3ePBV(NE9.7ICAH@CA\=5#+)Z6-
:eETUE/^4Y6?;b#?0S^WZ+bA>VTBJI/bZVNf4S>OaZ.P;cZ,@#9@#E-1NNb90955
61.WecR6D)6B(]QL0dL?I5B\Jdf9Z21QC+AUV8^E18+6JTT9,1)9Y<4<^PZcIU/:
V\I::0b:B_H<eLA+BQP,Q@H^WT=)T?M4G0297G]D@W^U:CT&GL7.SBc3-f\KK.]A
6HPBZdX1,1MD34D7UY:K()CG3)^ERN<,g]U6_34E==Y^UU\[(/;G5Cc_OQWb@-b<
L]+OaV2e,?3gcRc]6f9XcaR=e4G&(UGG,a6P(FR-P>325AB,7Y_f5bD4M7W8b86N
VNI@fI=&<Ge3+KJ_fT\PQ=<H;0ZFU>J9JL[0&8YD3D76FbNJY&,4OU+U/A,a5gbX
?TU#YZS[M/RTKE+TRJ<LY/QO(X@5=a;gFB1)9c<9HG\Dd/<IOaR@#P-eb=PKB;G3
b+EWKAJX,YRFATY.V,0Y-7CCf&X27#,4U/D9_)[K<ZW9@b;^::_CD0C@A-X]K3.G
131M[HFfQ9-6.4PK#\#9a,HU>HBB9W[[9?A<7[(bABNJM;D.cZ3-@CKGV1<E_KSB
bZ-DJP<X?,)3Y/BZN1dc_<aQ,EZY:ZgGD/91/UV4;D_^Tc,92e=G0+M+<=Rf/T&+
N[/](SbLJ4RY?4:CSXBQ:;>3HgDOE/N_3f-_M7b78;f+]>WaPK6NU.K_S[6O9ZQ^
[<aF+YSHdM^8KPJ91#H_XT&-V&+(XbKJ1588(HG5LP\H,1c#LHE1=:aD\Hg]I:C8
&/9<Be?#Oe<E@_Y0g/TELSJDR^RZX_S1?M9P+M=[X(a0SXDaV^&UI)GAK@\5-Y#J
XeFA=1AYNa[)e#>8&G&.7Y2W9=Afg9Sd:@]US-44Aa8Y9Y_+K\4U,5eaQ\^K-g,6
K+?ETYPP=AT.Ke4VcQ][C=K:=K-<81]PTb??Lc>72E7P-SG>gH6e/13Xg#_BCeUJ
#Z0WCF93#TMcHW,4[C.0#6fCF15BB/a6S:^SgJN^bE9:J-UK:D1E_R3XI$
`endprotected
endmodule

