//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2025 Fall
//   Lab01 Exercise		: Multi-Packet Channel Arbiter
//   Author     		: YU-CHEN CHANG
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : V1.0 (Release Date: 2025-09)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`define CYCLE_TIME 36.5

`ifdef RTL
	`define PATTERN_NUM 1
`endif
`ifdef GATE
	`define PATTERN_NUM 1
`endif

module PATTERN(
  // Output signals
    packets,
    channel_load,
    channel_capacity,
    KEY,
  // Input signals
    grant_channel 
);

//================================================================
//   INPUT AND OUTPUT DECLARATION                         
//================================================================
output reg [127:0] packets;
output reg  [11:0] channel_load;
output reg   [8:0] channel_capacity;
output reg  [63:0] KEY;

input [15:0] grant_channel ;

//================================================================
// parameters & integer
//================================================================
integer PATNUM = 1;
integer patcount;
integer input_file, output_file;
integer k,i,j;

//================================================================
// wire & registers 
//================================================================
reg [15:0] golden_packet [0:7];
reg [3:0] golden_channel_load[0:2];
reg [2:0] golden_channel_cap[0:2];

reg [1:0] golden_grant_channel[0:7];
reg [15:0] golden_grant_channel_a;
reg [63:0] golden_KEY;

//================================================================
// clock
//================================================================
reg clk;
real	CYCLE = `CYCLE_TIME;
always	#(CYCLE/2.0) clk = ~clk;
initial	clk = 0;

//================================================================
// Hint
//================================================================
// if you want to use c++/python to generate test data, here is 
// a sample format for you. You can change for your convinience.
/* 
input.txt format (using hex)
1. [PATTERN_NUM] 
repeat(PATTERN_NUM)
	1. [packet0]
    2. [packet1]
    3. [packet2]
    4. [packet3]
    5. [packet4]
    6. [packet5]
    7. [packet6]
    8. [packet7]
    9. [KEY]
    10.[channel_load0]
    11.[channel_load1]
    12.[channel_load2]
    13.[channel_capacity0]
    14.[channel_capacity1]
    15.[channel_capacity2]

 output.txt format (using hex or dec is ok, only range from 0~3)
 repeat(PATTERN_NUM)
    1. [grant_channel0]
    2. [grant_channel1]
    3. [grant_channel2]
    4. [grant_channel3]
    5. [grant_channel4]
    6. [grant_channel5]
    7. [grant_channel6]
    8. [grant_channel7]
*/

//================================================================
// initial
//================================================================
initial begin
    //please remember to save the original pattern
	input_file=$fopen("../00_TESTBED/input.txt","r");
    output_file=$fopen("../00_TESTBED/output.txt","r");

    packets = 'bx;
    channel_load = 'bx;

    repeat(5) @(negedge clk);

    k = $fscanf(input_file, "%d", PATNUM);

	for( patcount = 0; patcount < PATNUM; patcount++) begin		
        input_task;
        repeat(1) @(negedge clk);
		check_ans;
		// repeat($urandom_range(3, 5)) @(negedge clk);
        repeat(2) @(negedge clk);
        
	end
	display_pass;
    repeat(3) @(negedge clk);
    $finish;
end

//================================================================
// task
//================================================================

task input_task; begin
    for ( i = 0; i < 15; i++) begin
        if(i < 8)
        k = $fscanf(input_file, "%h", golden_packet[i]);
        else if(i < 9)
        k = $fscanf(input_file, "%h", golden_KEY);
        else if(i < 12)
        k = $fscanf(input_file, "%h", golden_channel_load[i-9]);
        else
        k = $fscanf(input_file, "%h", golden_channel_cap[i-12]);
    end
    

    packets = {golden_packet[7], golden_packet[6], golden_packet[5], golden_packet[4], 
               golden_packet[3], golden_packet[2], golden_packet[1], golden_packet[0]};
    
    KEY = golden_KEY;

    channel_load = {golden_channel_load[2], golden_channel_load[1], golden_channel_load[0]};

    channel_capacity = {golden_channel_cap[2], golden_channel_cap[1], golden_channel_cap[0]};

end endtask

task check_ans; begin
    for ( i = 0; i < 8; i++) begin
        k = $fscanf(output_file, "%h", golden_grant_channel[i]);
    end

    golden_grant_channel_a = {golden_grant_channel[7],golden_grant_channel[6], golden_grant_channel[5], golden_grant_channel[4],
                              golden_grant_channel[3],golden_grant_channel[2], golden_grant_channel[1], golden_grant_channel[0]};
    
    if (grant_channel !== golden_grant_channel_a) begin
        $display ("             \033[0;31mFAIL Pattern NO. %d\033[m         ", patcount);
        display_fail;
        $display ("   ------------------------------------------------------------------------");
        $display ("                                       FAIL                              ");
		$display("                                   PATTERN NO.%4d 	                      ", patcount);
        $display ("   Output should be : %b , your answer is : %b           ", golden_grant_channel_a, grant_channel);
        $display ("   ------------------------------------------------------------------------");
        #(200);
        $finish ;
    end
    else display_pass_gradient(patcount);
end endtask

task display_fail; begin
    $display("\n");
    $display("\n");
    
    $display("[38;2;54;61;67m█[0m[38;2;41;49;52m█[0m[38;2;40;48;51m█[0m[38;2;39;44;48m█[0m[38;2;34;41;47m█[0m[38;2;30;39;44m█[0m[38;2;41;46;50m█[0m[38;2;40;45;49m█[0m[38;2;43;48;52m█[0m[38;2;40;45;49m█[0m[38;2;39;44;48m█[0m[38;2;40;45;49m█[0m[38;2;46;51;55m█[0m[38;2;35;43;46m█[0m[38;2;42;50;53m█[0m[38;2;43;51;54m█[0m[38;2;44;52;55m█[0m[38;2;48;56;59m█[0m[38;2;41;49;52m█[0m[38;2;44;52;55m███[0m[38;2;39;47;50m██[0m[38;2;40;48;51m█[0m[38;2;42;47;51m█[0m[38;2;63;77;80m█[0m[38;2;36;44;47m█[0m[38;2;48;56;59m█[0m[38;2;47;55;58m█[0m[38;2;43;51;54m█[0m[38;2;42;50;53m█[0m[38;2;40;48;51m█[0m[38;2;36;41;45m█[0m[38;2;37;42;45m█[0m[38;2;48;56;59m█[0m[38;2;38;43;47m█[0m[38;2;37;42;46m█[0m[38;2;38;43;47m██[0m[38;2;41;46;50m█[0m[38;2;43;51;54m█[0m[38;2;46;51;55m█[0m[38;2;80;96;109m█[0m[38;2;50;58;60m█[0m[38;2;45;53;56m█[0m[38;2;46;54;57m█[0m[38;2;50;58;61m█[0m[38;2;39;44;48m██[0m[38;2;35;43;46m█[0m[38;2;43;51;54m█[0m[38;2;34;41;47m█[0m[38;2;37;42;46m██[0m[38;2;34;42;45m█[0m[38;2;74;87;95m█[0m[38;2;39;47;50m█[0m[38;2;39;44;48m█[0m[38;2;37;42;46m█[0m[38;2;41;46;50m█[0m[38;2;33;41;44m█[0m[38;2;49;57;60m█[0m[38;2;35;43;46m█[0m[38;2;39;44;48m█[0m[38;2;41;46;50m█[0m[38;2;47;55;58m█[0m[38;2;38;43;47m█[0m[38;2;41;46;50m█[0m[38;2;38;43;47m█[0m[38;2;44;49;53m█[0m[38;2;40;45;49m█[0m[38;2;38;46;49m█[0m[38;2;41;49;52m█[0m[38;2;39;47;50m██[0m[38;2;38;46;49m█[0m[38;2;51;59;62m█[0m[38;2;47;55;58m█[0m[38;2;46;54;57m███[0m[38;2;44;52;55m█[0m[38;2;53;61;64m█[0m[38;2;81;98;108m█[0m[38;2;45;53;56m█[0m[38;2;46;54;57m█[0m[38;2;51;59;62m█[0m[38;2;45;53;56m█[0m[38;2;43;51;54m█[0m[38;2;37;45;48m█[0m[38;2;41;49;52m█[0m[38;2;42;50;53m█[0m[38;2;46;54;57m█[0m[38;2;45;53;56m█[0m[38;2;50;58;61m█[0m[38;2;45;53;56m█[0m[38;2;46;54;57m█[0m[38;2;41;49;52m█[0m[38;2;48;56;59m█[0m");
$display("[38;2;50;58;61m█[0m[38;2;72;81;86m█[0m[38;2;51;59;62m█[0m[38;2;50;58;61m█[0m[38;2;51;59;62m█[0m[38;2;53;61;64m█[0m[38;2;94;107;115m█[0m[38;2;51;59;62m█[0m[38;2;50;58;61m█[0m[38;2;47;55;58m█[0m[38;2;46;54;57m█[0m[38;2;45;53;56m█[0m[38;2;47;55;58m█[0m[38;2;52;60;63m█[0m[38;2;72;80;83m█[0m[38;2;65;72;78m█[0m[38;2;71;79;82m█[0m[38;2;59;67;70m██[0m[38;2;58;66;69m█[0m[38;2;47;55;58m██[0m[38;2;50;58;61m█[0m[38;2;38;46;49m█[0m[38;2;34;42;45m█[0m[38;2;37;45;48m█[0m[38;2;41;49;52m█[0m[38;2;62;78;91m█[0m[38;2;37;42;46m█[0m[38;2;41;46;50m█[0m[38;2;37;42;46m█[0m[38;2;38;43;47m█[0m[38;2;36;41;45m█[0m[38;2;40;45;49m█[0m[38;2;38;43;47m█[0m[38;2;35;40;44m█[0m[38;2;37;44;50m█[0m[38;2;48;53;57m█[0m[38;2;46;51;55m█[0m[38;2;49;57;60m█[0m[38;2;45;53;56m██[0m[38;2;48;56;59m█[0m[38;2;51;56;60m█[0m[38;2;82;101;115m█[0m[38;2;50;58;61m██[0m[38;2;51;59;62m█[0m[38;2;47;55;58m█[0m[38;2;51;59;62m█[0m[38;2;49;57;60m█[0m[38;2;38;46;49m█[0m[38;2;39;47;50m█[0m[38;2;57;68;74m█[0m[38;2;42;50;53m█[0m[38;2;39;47;50m█[0m[38;2;36;44;47m█[0m[38;2;34;42;45m█[0m[38;2;40;45;49m█[0m[38;2;38;43;47m█[0m[38;2;39;44;48m█[0m[38;2;42;47;51m█[0m[38;2;47;52;56m█[0m[38;2;51;59;62m█[0m[38;2;38;46;49m█[0m[38;2;36;44;47m█[0m[38;2;40;48;51m█[0m[38;2;52;63;67m█[0m[38;2;46;51;55m█[0m[38;2;39;44;48m█[0m[38;2;38;46;49m█[0m[38;2;42;50;53m█[0m[38;2;39;47;50m█[0m[38;2;47;55;58m█[0m[38;2;48;56;59m█[0m[38;2;43;51;54m█[0m[38;2;40;48;51m█[0m[38;2;44;52;55m█[0m[38;2;48;56;59m█[0m[38;2;47;56;61m█[0m[38;2;49;57;60m█[0m[38;2;46;54;57m██[0m[38;2;47;55;58m█[0m[38;2;45;53;56m█[0m[38;2;99;112;120m█[0m[38;2;53;62;67m█[0m[38;2;43;51;54m█[0m[38;2;36;44;47m█[0m[38;2;38;43;47m█[0m[38;2;39;44;48m█[0m[38;2;35;40;44m█[0m[38;2;37;42;46m█[0m[38;2;36;41;45m█[0m[38;2;46;54;57m█[0m[38;2;44;52;55m█[0m[38;2;45;53;56m█[0m[38;2;46;54;57m█[0m[38;2;38;43;46m█[0m[38;2;37;42;45m█[0m");
$display("[38;2;50;58;61m█[0m[38;2;52;60;63m█[0m[38;2;50;61;65m█[0m[38;2;58;66;69m█[0m[38;2;53;61;64m█[0m[38;2;54;62;65m█[0m[38;2;47;57;59m█[0m[38;2;92;106;117m█[0m[38;2;51;59;62m███[0m[38;2;52;60;63m█[0m[38;2;51;59;62m█[0m[38;2;64;72;75m█[0m[38;2;72;82;84m█[0m[38;2;77;87;89m█[0m[38;2;68;77;82m█[0m[38;2;73;82;87m█[0m[38;2;65;74;79m█[0m[38;2;65;72;78m█[0m[38;2;45;53;56m█[0m[38;2;48;56;59m█[0m[38;2;45;53;56m█[0m[38;2;39;47;50m██[0m[38;2;41;49;52m█[0m[38;2;38;46;49m█[0m[38;2;35;43;46m█[0m[38;2;102;115;124m█[0m[38;2;38;43;47m██[0m[38;2;41;46;50m█[0m[38;2;37;42;46m█[0m[38;2;42;47;51m██[0m[38;2;36;41;45m█[0m[38;2;42;47;51m█[0m[38;2;33;44;46m█[0m[38;2;39;46;52m█[0m[38;2;44;52;55m█[0m[38;2;53;61;64m█[0m[38;2;46;54;57m█[0m[38;2;50;58;61m██[0m[38;2;50;54;57m█[0m[38;2;93;115;129m█[0m[38;2;50;55;59m█[0m[38;2;50;58;61m█[0m[38;2;51;59;62m█[0m[38;2;53;61;64m█[0m[38;2;49;57;60m█[0m[38;2;53;61;64m█[0m[38;2;50;58;61m█[0m[38;2;49;57;60m█[0m[38;2;84;101;111m█[0m[38;2;49;57;60m█[0m[38;2;37;45;48m█[0m[38;2;40;48;51m█[0m[38;2;39;47;50m█[0m[38;2;41;49;52m█[0m[38;2;38;46;49m█[0m[38;2;39;47;50m█[0m[38;2;43;48;52m█[0m[38;2;39;44;48m█[0m[38;2;42;50;53m██[0m[38;2;40;48;51m█[0m[38;2;44;52;54m█[0m[38;2;85;98;107m█[0m[38;2;52;59;65m█[0m[38;2;50;58;61m██[0m[38;2;51;59;62m█[0m[38;2;43;51;54m█[0m[38;2;48;56;59m█[0m[38;2;55;63;66m█[0m[38;2;48;56;59m█[0m[38;2;37;45;48m█[0m[38;2;38;46;49m█[0m[38;2;39;43;46m█[0m[38;2;69;80;86m█[0m[38;2;41;46;50m█[0m[38;2;40;45;49m█[0m[38;2;35;43;46m█[0m[38;2;34;42;44m█[0m[38;2;41;45;48m█[0m[38;2;15;24;29m█[0m[38;2;28;33;37m█[0m[38;2;36;41;45m██[0m[38;2;37;42;46m█[0m[38;2;39;44;48m█[0m[38;2;36;41;45m█[0m[38;2;37;42;46m█[0m[38;2;36;41;45m█[0m[38;2;41;45;48m█[0m[38;2;36;44;47m█[0m[38;2;35;43;46m█[0m[38;2;38;43;47m██[0m");
$display("[38;2;50;58;61m██[0m[38;2;52;60;63m█[0m[38;2;48;55;61m█[0m[38;2;60;69;76m█[0m[38;2;51;61;63m█[0m[38;2;55;63;66m█[0m[38;2;46;54;57m█[0m[38;2;74;92;104m█[0m[38;2;55;63;66m█[0m[38;2;47;55;58m█[0m[38;2;46;54;57m█[0m[38;2;70;78;81m█[0m[38;2;73;82;87m█[0m[38;2;63;73;75m█[0m[38;2;69;79;81m█[0m[38;2;60;70;72m█[0m[38;2;63;73;75m█[0m[38;2;67;77;79m█[0m[38;2;65;74;79m█[0m[38;2;62;70;73m█[0m[38;2;54;62;65m█[0m[38;2;46;51;55m█[0m[38;2;46;54;56m█[0m[38;2;38;46;48m█[0m[38;2;39;47;50m█[0m[38;2;33;41;44m█[0m[38;2;39;44;48m█[0m[38;2;40;45;49m█[0m[38;2;56;61;65m█[0m[38;2;36;40;43m█[0m[38;2;40;45;49m█[0m[38;2;37;42;46m█[0m[38;2;36;41;45m█[0m[38;2;44;49;53m█[0m[38;2;39;44;48m█[0m[38;2;41;46;50m█[0m[38;2;39;44;48m█[0m[38;2;36;41;45m█[0m[38;2;55;62;68m█[0m[38;2;37;42;48m█[0m[38;2;50;58;61m█[0m[38;2;54;62;65m█[0m[38;2;49;57;60m█[0m[38;2;47;55;58m█[0m[38;2;50;60;62m█[0m[38;2;98;111;120m█[0m[38;2;43;48;52m█[0m[38;2;46;54;57m█[0m[38;2;43;51;54m█[0m[38;2;47;55;58m█[0m[38;2;41;49;52m█[0m[38;2;48;56;59m█[0m[38;2;39;44;48m█[0m[38;2;44;49;53m█[0m[38;2;86;103;113m█[0m[38;2;47;52;55m█[0m[38;2;37;45;48m██[0m[38;2;37;42;46m█[0m[38;2;43;48;52m█[0m[38;2;38;43;47m█[0m[38;2;42;47;50m█[0m[38;2;53;61;64m█[0m[38;2;39;47;49m█[0m[38;2;55;62;68m█[0m[38;2;55;63;66m█[0m[38;2;48;56;59m█[0m[38;2;59;67;70m█[0m[38;2;98;108;118m█[0m[38;2;50;58;61m█[0m[38;2;51;60;65m█[0m[38;2;60;68;71m█[0m[38;2;45;53;56m█[0m[38;2;56;64;67m█[0m[38;2;54;62;65m█[0m[38;2;39;47;50m█[0m[38;2;37;45;48m█[0m[38;2;38;43;47m█[0m[38;2;36;41;45m█[0m[38;2;38;43;47m█[0m[38;2;72;86;95m█[0m[38;2;31;39;41m█[0m[38;2;43;48;52m█[0m[38;2;38;43;47m███[0m[38;2;34;44;46m█[0m[38;2;116;130;139m█[0m[38;2;39;47;50m█[0m[38;2;35;40;44m█[0m[38;2;49;54;58m█[0m[38;2;39;44;48m█[0m[38;2;37;42;46m█[0m[38;2;34;42;45m█[0m[38;2;43;51;54m█[0m[38;2;37;45;48m█[0m[38;2;39;47;50m█[0m[38;2;38;46;49m█[0m[38;2;45;53;56m█[0m");
$display("[38;2;46;54;57m█[0m[38;2;37;45;48m█[0m[38;2;44;52;55m█[0m[38;2;42;50;53m█[0m[38;2;41;49;52m█[0m[38;2;48;57;64m█[0m[38;2;49;57;60m██[0m[38;2;53;61;64m█[0m[38;2;72;85;93m█[0m[38;2;44;52;55m█[0m[38;2;52;60;63m█[0m[38;2;63;70;76m█[0m[38;2;75;84;89m█[0m[38;2;62;70;73m█[0m[38;2;64;72;75m█[0m[38;2;63;71;74m█[0m[38;2;56;64;67m█[0m[38;2;52;60;63m█[0m[38;2;61;70;75m█[0m[38;2;69;77;80m█[0m[38;2;62;70;73m██[0m[38;2;61;69;72m█[0m[38;2;41;50;55m█[0m[38;2;43;51;54m██[0m[38;2;36;44;47m█[0m[38;2;44;49;53m█[0m[38;2;35;40;44m█[0m[38;2;34;41;47m█[0m[38;2;31;39;42m█[0m[38;2;38;43;47m█[0m[38;2;37;42;46m█[0m[38;2;41;46;50m█[0m[38;2;36;41;45m█[0m[38;2;41;46;50m█[0m[38;2;36;44;47m█[0m[38;2;34;42;45m██[0m[38;2;36;44;46m█[0m[38;2;42;47;51m█[0m[38;2;40;45;49m█[0m[38;2;39;44;48m█[0m[38;2;43;48;52m█[0m[38;2;43;51;54m█[0m[38;2;39;47;50m██[0m[38;2;44;52;55m█[0m[38;2;45;53;56m█[0m[38;2;41;49;52m█[0m[38;2;40;48;51m█[0m[38;2;46;54;57m█[0m[38;2;33;41;44m█[0m[38;2;45;50;54m█[0m[38;2;41;49;52m█[0m[38;2;82;96;107m█[0m[38;2;45;53;56m█[0m[38;2;41;46;50m█[0m[38;2;37;45;48m█[0m[38;2;39;47;50m█[0m[38;2;41;49;52m█[0m[38;2;37;45;48m█[0m[38;2;51;59;62m█[0m[38;2;74;85;89m█[0m[38;2;52;59;65m█[0m[38;2;64;72;75m█[0m[38;2;48;56;59m█[0m[38;2;50;58;61m█[0m[38;2;56;64;67m█[0m[38;2;41;52;56m█[0m[38;2;48;56;59m█[0m[38;2;51;59;62m█[0m[38;2;48;56;59m█[0m[38;2;38;46;49m█[0m[38;2;39;47;50m██[0m[38;2;47;55;58m█[0m[38;2;41;46;50m██[0m[38;2;40;45;49m█[0m[38;2;39;44;47m█[0m[38;2;101;114;122m█[0m[38;2;44;49;52m█[0m[38;2;39;44;48m█[0m[38;2;37;42;46m█[0m[38;2;42;47;51m█[0m[38;2;36;45;50m█[0m[38;2;31;39;42m█[0m[38;2;87;104;114m█[0m[38;2;37;41;42m█[0m[38;2;36;41;45m█[0m[38;2;40;45;49m█[0m[38;2;41;46;50m█[0m[38;2;42;50;53m██[0m[38;2;43;51;54m██[0m[38;2;46;54;57m█[0m[38;2;45;53;56m█[0m");
$display("[38;2;41;49;52m█████[0m[38;2;33;41;43m█[0m[38;2;80;91;95m█[0m[38;2;45;50;54m█[0m[38;2;43;51;54m█[0m[38;2;50;58;61m█[0m[38;2;53;61;64m█[0m[38;2;67;77;79m█[0m[38;2;76;86;88m█[0m[38;2;65;75;77m█[0m[38;2;64;72;75m█[0m[38;2;65;73;76m█[0m[38;2;55;63;66m█[0m[38;2;63;73;75m█[0m[38;2;61;71;73m█[0m[38;2;61;69;72m██[0m[38;2;62;70;73m█[0m[38;2;54;62;65m█[0m[38;2;51;59;62m█[0m[38;2;50;58;61m█[0m[38;2;37;46;53m█[0m[38;2;52;61;66m█[0m[38;2;39;47;50m█[0m[38;2;40;48;51m█[0m[38;2;35;43;46m█[0m[38;2;34;39;43m█[0m[38;2;37;42;46m█[0m[38;2;42;47;51m█[0m[38;2;33;38;42m█[0m[38;2;41;46;50m█[0m[38;2;39;44;48m█[0m[38;2;36;41;45m█[0m[38;2;38;46;49m█[0m[38;2;39;47;50m█[0m[38;2;35;44;49m█[0m[38;2;41;48;56m█[0m[38;2;41;49;52m█[0m[38;2;47;55;58m█[0m[38;2;37;45;48m█[0m[38;2;36;41;45m█[0m[38;2;43;51;54m█[0m[38;2;40;48;51m█[0m[38;2;42;50;53m█[0m[38;2;36;44;47m█[0m[38;2;40;48;51m█[0m[38;2;44;49;53m█[0m[38;2;41;46;50m█[0m[38;2;37;45;48m█[0m[38;2;45;53;56m█[0m[38;2;37;44;50m█[0m[38;2;40;48;51m█[0m[38;2;41;49;52m█[0m[38;2;43;52;57m█[0m[38;2;39;47;50m██[0m[38;2;38;46;49m█[0m[38;2;37;45;48m█[0m[38;2;43;51;54m█[0m[38;2;44;52;55m█[0m[38;2;53;61;64m█[0m[38;2;45;54;61m█[0m[38;2;51;59;62m█[0m[38;2;43;51;54m█[0m[38;2;48;56;59m█[0m[38;2;50;58;61m█[0m[38;2;41;49;52m█[0m[38;2;23;36;42m█[0m[38;2;29;40;42m█[0m[38;2;44;52;55m█[0m[38;2;47;55;58m█[0m[38;2;41;49;52m██[0m[38;2;36;44;47m█[0m[38;2;40;45;49m█[0m[38;2;45;50;54m█[0m[38;2;37;42;46m█[0m[38;2;43;48;52m█[0m[38;2;44;49;53m█[0m[38;2;95;105;115m█[0m[38;2;39;49;51m█[0m[38;2;38;46;49m█[0m[38;2;40;45;49m█[0m[38;2;46;51;55m█[0m[38;2;38;43;47m█[0m[38;2;42;47;51m█[0m[38;2;94;112;122m█[0m[38;2;41;46;49m█[0m[38;2;39;47;50m█[0m[38;2;37;45;48m█[0m[38;2;43;51;54m█[0m[38;2;39;47;49m█[0m[38;2;53;60;66m█[0m[38;2;40;48;51m█[0m[38;2;39;47;50m█[0m[38;2;45;53;56m█[0m");
$display("[38;2;46;56;58m█[0m[38;2;55;63;66m█[0m[38;2;51;59;62m█[0m[38;2;44;52;55m█[0m[38;2;41;49;52m█[0m[38;2;43;51;54m█[0m[38;2;48;56;58m█[0m[38;2;76;86;95m█[0m[38;2;61;70;75m█[0m[38;2;62;72;74m██[0m[38;2;66;76;78m█[0m[38;2;60;70;72m█[0m[38;2;65;73;76m█[0m[38;2;62;70;73m█[0m[38;2;63;71;74m█[0m[38;2;59;67;70m█[0m[38;2;59;69;71m█[0m[38;2;66;76;78m█[0m[38;2;58;66;69m█[0m[38;2;57;65;68m█[0m[38;2;54;62;65m█[0m[38;2;52;60;63m█[0m[38;2;56;64;67m█[0m[38;2;51;59;62m█[0m[38;2;51;58;64m█[0m[38;2;56;64;67m█[0m[38;2;65;78;86m█[0m[38;2;50;58;61m█[0m[38;2;44;52;55m█[0m[38;2;45;53;56m█[0m[38;2;43;51;54m█[0m[38;2;39;47;50m█[0m[38;2;47;55;58m█[0m[38;2;64;74;76m█[0m[38;2;43;51;54m█[0m[38;2;39;47;50m█[0m[38;2;50;58;61m█[0m[38;2;48;56;59m█[0m[38;2;53;61;64m█[0m[38;2;53;62;67m█[0m[38;2;98;112;121m█[0m[38;2;58;66;69m█[0m[38;2;60;68;71m█[0m[38;2;55;63;66m█[0m[38;2;50;58;61m█[0m[38;2;35;43;46m█[0m[38;2;43;51;54m██[0m[38;2;39;47;50m██[0m[38;2;40;48;51m█[0m[38;2;44;52;55m██[0m[38;2;50;58;61m█[0m[38;2;37;46;53m█[0m[38;2;44;52;55m█[0m[38;2;43;51;54m█[0m[38;2;40;48;51m██[0m[38;2;47;55;58m█[0m[38;2;55;63;66m█[0m[38;2;52;60;63m█[0m[38;2;53;61;64m█[0m[38;2;56;64;67m█[0m[38;2;52;60;63m█[0m[38;2;61;70;75m█[0m[38;2;49;60;66m█[0m[38;2;52;61;66m█[0m[38;2;57;65;68m█[0m[38;2;55;63;66m█[0m[38;2;53;61;64m█[0m[38;2;53;63;65m█[0m[38;2;112;127;134m█[0m[38;2;51;56;59m█[0m[38;2;43;51;54m█[0m[38;2;48;56;59m█[0m[38;2;47;55;58m█[0m[38;2;40;48;51m█[0m[38;2;47;55;58m█[0m[38;2;40;48;51m█[0m[38;2;44;52;55m█[0m[38;2;45;53;56m█[0m[38;2;43;51;54m█[0m[38;2;29;42;48m█[0m[38;2;45;56;62m█[0m[38;2;39;44;48m█[0m[38;2;42;50;53m█[0m[38;2;41;49;52m█[0m[38;2;36;41;45m█[0m[38;2;41;46;50m█[0m[38;2;39;47;50m██[0m[38;2;42;50;53m█[0m[38;2;40;48;51m█[0m[38;2;37;45;48m█[0m[38;2;41;49;52m█[0m[38;2;41;48;54m█[0m[38;2;38;46;49m██[0m");
$display("[38;2;62;70;73m█[0m[38;2;68;78;87m█[0m[38;2;62;70;73m█[0m[38;2;64;72;75m█[0m[38;2;60;68;71m█[0m[38;2;59;69;71m█[0m[38;2;57;65;68m█[0m[38;2;64;72;75m█[0m[38;2;99;113;124m█[0m[38;2;69;77;80m█[0m[38;2;59;67;70m█[0m[38;2;65;73;76m█[0m[38;2;64;72;75m█[0m[38;2;61;69;72m█[0m[38;2;56;64;67m█[0m[38;2;62;70;73m█[0m[38;2;65;73;76m█[0m[38;2;58;66;69m█[0m[38;2;62;70;73m█[0m[38;2;61;69;72m█[0m[38;2;62;70;73m█[0m[38;2;54;62;65m█[0m[38;2;59;67;70m█[0m[38;2;54;62;65m█[0m[38;2;53;61;64m█[0m[38;2;46;54;57m█[0m[38;2;58;66;69m█[0m[38;2;58;68;70m█[0m[38;2;84;101;111m█[0m[38;2;49;58;63m█[0m[38;2;53;61;64m█[0m[38;2;54;62;65m█[0m[38;2;46;54;57m█[0m[38;2;48;56;59m█[0m[38;2;44;52;55m█[0m[38;2;46;54;57m█[0m[38;2;56;66;68m█[0m[38;2;47;55;58m█[0m[38;2;44;52;55m█[0m[38;2;50;58;61m█[0m[38;2;55;63;66m█[0m[38;2;62;72;74m█[0m[38;2;90;107;117m█[0m[38;2;65;75;77m█[0m[38;2;55;63;66m█[0m[38;2;54;62;65m██[0m[38;2;51;59;62m█[0m[38;2;52;60;63m█[0m[38;2;60;68;71m█[0m[38;2;60;69;74m█[0m[38;2;58;69;75m█[0m[38;2;55;63;66m█[0m[38;2;51;59;62m█[0m[38;2;45;53;56m█[0m[38;2;49;56;62m█[0m[38;2;71;84;92m█[0m[38;2;50;58;61m█[0m[38;2;54;62;65m█[0m[38;2;53;61;64m█[0m[38;2;51;59;62m█[0m[38;2;55;63;66m█[0m[38;2;51;59;62m██[0m[38;2;64;72;75m█[0m[38;2;55;63;66m█[0m[38;2;57;65;68m█[0m[38;2;60;69;74m█[0m[38;2;87;100;108m█[0m[38;2;54;62;65m█[0m[38;2;58;66;69m█[0m[38;2;53;61;64m█[0m[38;2;51;61;63m█[0m[38;2;57;67;69m█[0m[38;2;93;110;120m█[0m[38;2;61;69;72m██[0m[38;2;62;70;73m█[0m[38;2;57;65;68m█[0m[38;2;60;68;71m██[0m[38;2;52;60;63m█[0m[38;2;46;54;57m█[0m[38;2;39;47;50m█[0m[38;2;43;53;55m█[0m[38;2;48;58;60m█[0m[38;2;85;98;107m█[0m[38;2;43;51;54m█[0m[38;2;60;68;71m█[0m[38;2;54;62;65m█[0m[38;2;48;56;59m█[0m[38;2;42;50;53m█[0m[38;2;41;49;52m█[0m[38;2;42;50;53m█[0m[38;2;43;51;54m█[0m[38;2;41;49;52m█[0m[38;2;43;51;54m██[0m[38;2;64;71;77m█[0m[38;2;52;63;67m█[0m");
$display("[38;2;62;70;73m█[0m[38;2;63;71;74m█[0m[38;2;89;102;110m█[0m[38;2;61;69;72m█[0m[38;2;59;67;70m█[0m[38;2;62;70;73m█[0m[38;2;65;73;76m█[0m[38;2;62;70;73m█[0m[38;2;63;71;74m█[0m[38;2;97;115;129m█[0m[38;2;62;69;75m█[0m[38;2;61;69;72m█[0m[38;2;62;70;73m█[0m[38;2;58;66;69m█[0m[38;2;63;71;74m█[0m[38;2;62;70;73m█[0m[38;2;66;74;77m█[0m[38;2;62;72;74m█[0m[38;2;57;67;69m█[0m[38;2;55;63;66m█[0m[38;2;53;61;64m█[0m[38;2;58;66;69m█[0m[38;2;57;65;68m█[0m[38;2;58;66;69m█[0m[38;2;55;63;66m█[0m[38;2;64;72;75m█[0m[38;2;59;67;70m█[0m[38;2;71;79;82m█[0m[38;2;64;71;77m█[0m[38;2;75;94;109m█[0m[38;2;52;60;63m█[0m[38;2;53;61;64m█[0m[38;2;54;62;65m█[0m[38;2;47;55;58m█[0m[38;2;51;59;62m█[0m[38;2;52;60;63m█[0m[38;2;57;65;68m█[0m[38;2;77;86;93m█[0m[38;2;65;74;79m█[0m[38;2;60;68;71m█[0m[38;2;61;69;72m█[0m[38;2;74;81;87m█[0m[38;2;62;73;77m█[0m[38;2;116;132;145m█[0m[38;2;60;68;71m█[0m[38;2;65;73;76m█[0m[38;2;60;68;71m█[0m[38;2;65;73;76m█[0m[38;2;64;72;75m█[0m[38;2;60;68;71m█[0m[38;2;61;71;73m█[0m[38;2;59;70;74m█[0m[38;2;64;73;78m█[0m[38;2;65;73;76m█[0m[38;2;70;78;81m█[0m[38;2;61;71;73m█[0m[38;2;61;73;73m█[0m[38;2;89;102;108m█[0m[38;2;68;76;79m█[0m[38;2;62;72;74m█[0m[38;2;58;68;70m█[0m[38;2;50;58;61m█[0m[38;2;51;59;62m█[0m[38;2;60;68;71m█[0m[38;2;53;61;64m█[0m[38;2;56;64;67m█[0m[38;2;54;62;65m█[0m[38;2;52;60;63m█[0m[38;2;58;66;69m█[0m[38;2;84;99;106m█[0m[38;2;58;66;69m██[0m[38;2;56;64;67m█[0m[38;2;58;69;75m█[0m[38;2;69;77;80m█[0m[38;2;99;113;122m█[0m[38;2;58;68;70m█[0m[38;2;60;68;71m█[0m[38;2;62;70;73m█[0m[38;2;59;67;70m█[0m[38;2;60;68;71m█[0m[38;2;58;66;69m█[0m[38;2;67;75;78m█[0m[38;2;54;62;65m█[0m[38;2;57;65;68m█[0m[38;2;59;67;70m█[0m[38;2;52;61;66m█[0m[38;2;99;116;126m█[0m[38;2;65;73;75m█[0m[38;2;61;69;72m█[0m[38;2;65;73;76m█[0m[38;2;64;74;76m█[0m[38;2;59;67;70m█[0m[38;2;57;65;68m█[0m[38;2;55;63;66m█[0m[38;2;54;62;65m█[0m[38;2;56;64;67m██[0m[38;2;48;56;59m█[0m[38;2;57;65;68m█[0m");
$display("[38;2;59;69;71m█[0m[38;2;61;71;73m██[0m[38;2;96;115;122m█[0m[38;2;61;72;76m█[0m[38;2;61;69;72m██[0m[38;2;62;70;73m██[0m[38;2;64;75;81m█[0m[38;2;67;80;86m█[0m[38;2;55;65;67m█[0m[38;2;59;68;75m█[0m[38;2;62;72;74m█[0m[38;2;57;67;69m█[0m[38;2;67;77;79m█[0m[38;2;56;66;68m█[0m[38;2;67;80;86m█[0m[38;2;66;75;82m█[0m[38;2;68;77;82m█[0m[38;2;61;71;72m█[0m[38;2;64;75;79m█[0m[38;2;62;72;74m█[0m[38;2;61;71;73m█[0m[38;2;66;76;78m█[0m[38;2;65;74;79m█[0m[38;2;72;81;86m█[0m[38;2;66;75;80m█[0m[38;2;60;69;74m█[0m[38;2;70;79;84m█[0m[38;2;109;127;141m█[0m[38;2;65;75;77m█[0m[38;2;71;82;86m█[0m[38;2;72;81;86m█[0m[38;2;70;79;84m█[0m[38;2;79;88;93m█[0m[38;2;66;75;80m█[0m[38;2;65;75;76m█[0m[38;2;63;74;80m█[0m[38;2;69;76;82m█[0m[38;2;59;69;78m█[0m[38;2;66;74;77m█[0m[38;2;63;72;77m█[0m[38;2;77;86;91m█[0m[38;2;86;103;110m█[0m[38;2;59;69;71m█[0m[38;2;58;68;70m█[0m[38;2;59;68;73m█[0m[38;2;67;77;79m█[0m[38;2;60;70;72m█[0m[38;2;65;76;78m█[0m[38;2;63;73;75m█[0m[38;2;70;80;82m█[0m[38;2;59;72;78m█[0m[38;2;77;84;90m█[0m[38;2;25;16;9m█[0m[38;2;44;32;20m█[0m[38;2;34;22;10m█[0m[38;2;14;11;4m█[0m[38;2;70;83;89m█[0m[38;2;71;78;84m█[0m[38;2;73;82;87m█[0m[38;2;66;75;80m█[0m[38;2;70;79;84m█[0m[38;2;52;61;66m█[0m[38;2;51;61;63m█[0m[38;2;57;67;69m█[0m[38;2;57;65;68m█[0m[38;2;55;63;66m█[0m[38;2;57;67;69m█[0m[38;2;88;101;110m█[0m[38;2;64;71;77m█[0m[38;2;64;72;75m█[0m[38;2;70;78;81m█[0m[38;2;54;62;65m█[0m[38;2;59;69;70m█[0m[38;2;102;116;129m█[0m[38;2;54;64;66m█[0m[38;2;61;69;72m█[0m[38;2;57;65;68m██[0m[38;2;61;69;72m█[0m[38;2;55;62;68m█[0m[38;2;58;66;69m██[0m[38;2;57;65;68m█[0m[38;2;53;61;64m█[0m[38;2;57;65;68m█[0m[38;2;111;129;141m█[0m[38;2;65;75;77m█[0m[38;2;58;65;71m█[0m[38;2;60;68;71m█[0m[38;2;56;66;68m█[0m[38;2;72;83;87m█[0m[38;2;53;61;64m█[0m[38;2;54;62;65m█[0m[38;2;57;65;68m█[0m[38;2;55;63;66m█[0m[38;2;59;69;71m█[0m[38;2;68;78;80m█[0m");
$display("[38;2;61;70;75m█[0m[38;2;65;74;79m█[0m[38;2;56;66;68m█[0m[38;2;58;68;70m█[0m[38;2;99;113;124m█[0m[38;2;65;73;76m█[0m[38;2;66;74;77m█[0m[38;2;62;70;73m█[0m[38;2;73;81;84m█[0m[38;2;58;66;69m█[0m[38;2;62;70;73m█[0m[38;2;58;69;75m█[0m[38;2;57;68;72m█[0m[38;2;55;65;67m█[0m[38;2;58;68;70m██[0m[38;2;70;79;84m█[0m[38;2;23;16;8m█[0m[38;2;36;22;9m█[0m[38;2;34;22;10m█[0m[38;2;38;26;14m█[0m[38;2;36;24;12m█[0m[38;2;33;21;7m█[0m[38;2;12;9;4m█[0m[38;2;75;86;92m█[0m[38;2;79;86;94m█[0m[38;2;78;90;88m█[0m[38;2;74;83;88m█[0m[38;2;76;85;90m█[0m[38;2;71;80;85m█[0m[38;2;79;88;93m█[0m[38;2;89;103;112m█[0m[38;2;72;79;85m█[0m[38;2;74;83;88m█[0m[38;2;62;71;76m█[0m[38;2;70;79;84m█[0m[38;2;67;76;81m█[0m[38;2;77;86;91m█[0m[38;2;68;77;82m█[0m[38;2;67;76;81m█[0m[38;2;91;104;112m█[0m[38;2;66;76;78m█[0m[38;2;68;77;82m█[0m[38;2;66;75;80m█[0m[38;2;63;72;77m█[0m[38;2;68;77;82m█[0m[38;2;69;78;83m█[0m[38;2;72;83;85m█[0m[38;2;69;72;79m█[0m[38;2;75;84;83m█[0m[38;2;39;27;15m█[0m[38;2;36;22;9m█[0m[38;2;36;22;11m█[0m[38;2;34;25;8m█[0m[38;2;37;24;15m█[0m[38;2;17;0;0m█[0m[38;2;200;169;123m█[0m[38;2;77;48;16m█[0m[38;2;28;23;3m█[0m[38;2;33;23;13m█[0m[38;2;34;25;18m█[0m[38;2;80;87;97m█[0m[38;2;72;81;86m█[0m[38;2;67;76;81m█[0m[38;2;69;80;84m█[0m[38;2;97;111;120m█[0m[38;2;68;77;82m██[0m[38;2;67;76;81m█[0m[38;2;64;73;78m█[0m[38;2;69;77;80m█[0m[38;2;83;96;104m█[0m[38;2;62;71;76m█[0m[38;2;61;70;75m█[0m[38;2;60;69;74m█[0m[38;2;62;71;76m█[0m[38;2;60;69;74m█[0m[38;2;59;69;71m█[0m[38;2;66;76;78m█[0m[38;2;58;68;70m█[0m[38;2;56;64;67m█[0m[38;2;58;66;69m█[0m[38;2;57;65;68m█[0m[38;2;56;66;68m█[0m[38;2;57;65;68m█[0m[38;2;59;67;70m█[0m[38;2;53;61;64m█[0m[38;2;56;66;68m█[0m[38;2;65;75;77m█[0m[38;2;98;115;125m█[0m[38;2;57;67;69m█[0m[38;2;66;74;77m█[0m[38;2;54;62;65m█[0m[38;2;55;63;66m█[0m[38;2;81;91;100m█[0m[38;2;57;64;70m█[0m[38;2;62;69;75m█[0m[38;2;58;68;70m█[0m[38;2;71;80;85m█[0m[38;2;67;76;81m█[0m");
$display("[38;2;77;86;91m█[0m[38;2;74;83;88m█[0m[38;2;66;75;80m█[0m[38;2;64;74;76m██[0m[38;2;94;108;119m█[0m[38;2;48;61;67m█[0m[38;2;62;72;74m█[0m[38;2;60;68;71m█[0m[38;2;74;82;85m█[0m[38;2;60;68;71m█[0m[38;2;64;74;76m█[0m[38;2;65;75;77m█[0m[38;2;66;76;78m█[0m[38;2;67;76;81m█[0m[38;2;81;90;95m█[0m[38;2;32;25;17m█[0m[38;2;36;23;14m█[0m[38;2;24;2;0m█[0m[38;2;172;130;70m█[0m[38;2;183;142;78m█[0m[38;2;190;148;90m█[0m[38;2;189;156;113m█[0m[38;2;29;27;2m█[0m[38;2;37;19;17m█[0m[38;2;35;23;11m█[0m[38;2;34;21;12m█[0m[38;2;45;33;21m█[0m[38;2;97;102;105m█[0m[38;2;71;80;85m█[0m[38;2;76;87;91m█[0m[38;2;70;79;84m██[0m[38;2;80;89;94m█[0m[38;2;89;94;98m█[0m[38;2;76;90;93m█[0m[38;2;87;101;104m█[0m[38;2;81;94;100m█[0m[38;2;68;79;85m█[0m[38;2;73;88;93m█[0m[38;2;77;92;97m█[0m[38;2;72;87;92m█[0m[38;2;81;96;99m█[0m[38;2;68;86;90m█[0m[38;2;74;85;89m█[0m[38;2;69;78;77m█[0m[38;2;60;73;79m█[0m[38;2;34;22;10m█[0m[38;2;35;29;17m█[0m[38;2;39;22;12m█[0m[38;2;29;16;26m█[0m[38;2;192;142;89m█[0m[38;2;183;143;84m█[0m[38;2;181;139;81m█[0m[38;2;185;143;85m█[0m[38;2;183;143;84m█[0m[38;2;183;141;83m█[0m[38;2;186;144;86m█[0m[38;2;174;129;74m█[0m[38;2;34;25;18m█[0m[38;2;36;24;10m█[0m[38;2;31;31;29m█[0m[38;2;88;99;103m█[0m[38;2;85;96;100m█[0m[38;2;72;82;84m█[0m[38;2;66;77;83m█[0m[38;2;105;122;132m█[0m[38;2;70;79;84m██[0m[38;2;69;78;83m█[0m[38;2;70;79;84m█[0m[38;2;85;94;99m█[0m[38;2;81;92;98m█[0m[38;2;72;81;86m█[0m[38;2;75;84;89m█[0m[38;2;74;83;88m██[0m[38;2;73;82;87m█[0m[38;2;77;86;91m█[0m[38;2;71;80;85m█[0m[38;2;74;83;88m█[0m[38;2;64;74;76m█[0m[38;2;61;71;73m█[0m[38;2;60;70;72m█[0m[38;2;77;87;96m█[0m[38;2;65;75;77m█[0m[38;2;64;74;76m██[0m[38;2;58;68;70m█[0m[38;2;56;66;68m█[0m[38;2;63;73;75m█[0m[38;2;61;69;72m█[0m[38;2;69;77;80m█[0m[38;2;62;70;73m█[0m[38;2;62;72;74m█[0m[38;2;57;70;76m█[0m[38;2;63;72;77m█[0m[38;2;69;78;83m█[0m[38;2;68;77;82m█[0m[38;2;69;78;83m█[0m");
$display("[38;2;81;90;95m█[0m[38;2;78;87;92m█[0m[38;2;76;87;91m█[0m[38;2;80;89;94m█[0m[38;2;79;88;93m█[0m[38;2;78;87;92m█[0m[38;2;78;89;95m█[0m[38;2;69;82;90m█[0m[38;2;62;71;76m█[0m[38;2;58;67;72m█[0m[38;2;78;87;92m█[0m[38;2;69;78;83m█[0m[38;2;89;98;103m█[0m[38;2;84;93;98m█[0m[38;2;82;91;96m██[0m[38;2;34;20;7m█[0m[38;2;31;23;2m█[0m[38;2;179;133;83m█[0m[38;2;180;139;85m█[0m[38;2;174;133;77m█[0m[38;2;179;138;82m█[0m[38;2;184;144;85m█[0m[38;2;188;148;89m█[0m[38;2;174;134;75m█[0m[38;2;181;140;84m█[0m[38;2;182;135;79m█[0m[38;2;14;0;0m█[0m[38;2;32;21;17m█[0m[38;2;32;23;8m█[0m[38;2;32;22;10m█[0m[38;2;38;26;14m█[0m[38;2;37;20;10m█[0m[38;2;37;25;13m█[0m[38;2;34;22;10m██[0m[38;2;39;27;15m█[0m[38;2;31;22;7m█[0m[38;2;33;23;14m█[0m[38;2;37;18;11m█[0m[38;2;44;23;18m█[0m[38;2;40;21;15m█[0m[38;2;41;27;18m█[0m[38;2;35;22;6m█[0m[38;2;35;23;11m███[0m[38;2;36;22;13m█[0m[38;2;181;141;80m█[0m[38;2;183;140;85m█[0m[38;2;181;139;81m█[0m[38;2;186;144;86m██[0m[38;2;187;146;92m█[0m[38;2;185;146;89m█[0m[38;2;26;17;10m█[0m[38;2;196;166;114m█[0m[38;2;182;136;84m█[0m[38;2;185;143;85m█[0m[38;2;193;149;86m█[0m[38;2;35;28;12m█[0m[38;2;35;23;11m█[0m[38;2;85;96;100m█[0m[38;2;90;101;105m██[0m[38;2;85;96;100m█[0m[38;2;75;88;96m█[0m[38;2;110;127;137m█[0m[38;2;75;86;90m█[0m[38;2;88;99;103m█[0m[38;2;89;100;104m█[0m[38;2;85;94;99m█[0m[38;2;78;89;93m█[0m[38;2;81;92;96m██[0m[38;2;84;93;98m█[0m[38;2;83;92;97m█[0m[38;2;84;95;99m█[0m[38;2;88;99;103m█[0m[38;2;85;96;100m█[0m[38;2;84;93;98m█[0m[38;2;89;98;103m█[0m[38;2;86;95;100m██[0m[38;2;85;94;99m█[0m[38;2;101;115;124m█[0m[38;2;76;85;90m█[0m[38;2;66;75;80m█[0m[38;2;63;72;77m█[0m[38;2;66;76;78m█[0m[38;2;60;70;72m█[0m[38;2;58;66;69m█[0m[38;2;61;71;73m█[0m[38;2;60;70;72m█[0m[38;2;69;79;81m█[0m[38;2;64;71;77m█[0m[38;2;53;64;70m█[0m[38;2;81;90;95m█[0m[38;2;76;85;90m█[0m[38;2;69;78;83m█[0m");
$display("[38;2;86;95;100m█[0m[38;2;80;89;94m█[0m[38;2;86;95;100m█[0m[38;2;78;89;93m█[0m[38;2;80;91;95m█[0m[38;2;83;92;97m█[0m[38;2;79;90;92m█[0m[38;2;64;77;83m█[0m[38;2;106;123;131m█[0m[38;2;74;83;88m█[0m[38;2;78;87;92m█[0m[38;2;80;89;94m█[0m[38;2;85;94;99m█[0m[38;2;81;90;95m█[0m[38;2;80;91;95m█[0m[38;2;68;79;85m█[0m[38;2;36;24;12m█[0m[38;2;36;23;17m█[0m[38;2;169;126;75m█[0m[38;2;166;125;71m█[0m[38;2;40;26;25m█[0m[38;2;209;178;121m█[0m[38;2;185;145;86m█[0m[38;2;179;138;82m█[0m[38;2;188;147;91m█[0m[38;2;181;139;81m█[0m[38;2;176;134;76m█[0m[38;2;179;140;73m█[0m[38;2;35;22;14m█[0m[38;2;30;27;10m█[0m[38;2;45;30;23m█[0m[38;2;218;180;131m█[0m[38;2;181;145;83m█[0m[38;2;177;139;77m█[0m[38;2;182;131;78m█[0m[38;2;188;149;84m█[0m[38;2;180;144;84m█[0m[38;2;182;142;83m█[0m[38;2;179;139;80m█[0m[38;2;180;140;81m██[0m[38;2;186;144;86m█[0m[38;2;187;147;88m█[0m[38;2;191;146;87m█[0m[38;2;37;24;7m█[0m[38;2;21;5;0m█[0m[38;2;182;137;82m█[0m[38;2;182;142;83m█[0m[38;2;191;149;91m█[0m[38;2;182;140;82m█[0m[38;2;182;142;83m█[0m[38;2;184;144;85m█[0m[38;2;187;137;76m█[0m[38;2;38;25;8m█[0m[38;2;35;20;13m█[0m[38;2;111;139;151m█[0m[38;2;120;138;148m█[0m[38;2;182;137;78m█[0m[38;2;182;140;82m█[0m[38;2;183;143;84m█[0m[38;2;35;27;24m█[0m[38;2;28;20;7m█[0m[38;2;92;103;107m██[0m[38;2;90;101;105m█[0m[38;2;87;98;102m█[0m[38;2;92;101;106m█[0m[38;2;88;99;103m█[0m[38;2;86;97;101m█[0m[38;2;81;92;96m█[0m[38;2;76;91;94m█[0m[38;2;14;11;4m█[0m[38;2;38;24;13m█[0m[38;2;37;25;13m██[0m[38;2;38;26;14m█[0m[38;2;31;19;7m█[0m[38;2;37;25;13m█[0m[38;2;35;25;13m█[0m[38;2;39;27;15m█[0m[38;2;43;29;16m█[0m[38;2;32;25;15m█[0m[38;2;98;108;110m█[0m[38;2;87;98;102m█[0m[38;2;84;95;99m█[0m[38;2;87;96;101m█[0m[38;2;101;115;118m█[0m[38;2;88;97;102m█[0m[38;2;84;93;98m█[0m[38;2;65;74;79m█[0m[38;2;83;92;99m█[0m[38;2;65;74;79m█[0m[38;2;70;78;81m█[0m[38;2;75;83;86m█[0m[38;2;83;92;97m█[0m[38;2;62;71;76m█[0m[38;2;89;98;103m█[0m[38;2;82;93;99m█[0m[38;2;86;97;101m█[0m[38;2;84;95;99m█[0m");
$display("[38;2;108;121;127m█[0m[38;2;91;100;105m█[0m[38;2;78;89;93m█[0m[38;2;82;93;97m█[0m[38;2;73;84;88m█[0m[38;2;73;82;87m█[0m[38;2;72;81;86m█[0m[38;2;73;82;87m█[0m[38;2;65;78;86m█[0m[38;2;113;129;142m█[0m[38;2;75;85;87m█[0m[38;2;75;84;89m█[0m[38;2;74;83;88m█[0m[38;2;82;91;96m█[0m[38;2;81;90;95m█[0m[38;2;93;106;112m█[0m[38;2;34;22;10m█[0m[38;2;14;8;0m█[0m[38;2;153;109;60m█[0m[38;2;165;125;74m█[0m[38;2;161;117;70m█[0m[38;2;30;23;4m█[0m[38;2;37;24;16m█[0m[38;2;184;144;85m█[0m[38;2;186;146;87m█[0m[38;2;184;142;84m█[0m[38;2;177;135;77m█[0m[38;2;187;146;90m█[0m[38;2;184;141;86m█[0m[38;2;185;147;85m█[0m[38;2;185;145;86m█[0m[38;2;179;137;79m█[0m[38;2;183;141;83m█[0m[38;2;179;139;80m█[0m[38;2;187;148;89m█[0m[38;2;181;142;83m█[0m[38;2;182;141;85m█[0m[38;2;183;141;83m█[0m[38;2;189;147;89m█[0m[38;2;185;145;86m█[0m[38;2;188;148;89m█[0m[38;2;193;153;94m█[0m[38;2;189;149;90m█[0m[38;2;183;143;84m█[0m[38;2;192;152;91m█[0m[38;2;182;142;83m█[0m[38;2;175;135;76m█[0m[38;2;185;143;85m█[0m[38;2;180;140;81m█[0m[38;2;183;143;84m█[0m[38;2;183;141;83m█[0m[38;2;195;152;97m█[0m[38;2;34;26;13m█[0m[38;2;36;18;4m█[0m[38;2;112;126;139m█[0m[38;2;115;135;146m█[0m[38;2;119;138;152m█[0m[38;2;182;137;80m█[0m[38;2;179;137;79m█[0m[38;2;181;141;80m█[0m[38;2;206;174;115m█[0m[38;2;38;26;14m█[0m[38;2;29;18;14m█[0m[38;2;100;103;110m█[0m[38;2;87;98;102m█[0m[38;2;88;99;103m█[0m[38;2;97;108;112m█[0m[38;2;96;107;113m█[0m[38;2;87;98;104m█[0m[38;2;42;26;10m█[0m[38;2;33;25;12m█[0m[38;2;34;24;14m█[0m[38;2;171;133;70m█[0m[38;2;182;141;87m█[0m[38;2;183;145;83m█[0m[38;2;182;144;81m█[0m[38;2;180;140;89m█[0m[38;2;180;141;82m█[0m[38;2;184;142;82m█[0m[38;2;183;137;85m█[0m[38;2;189;144;89m█[0m[38;2;21;0;0m█[0m[38;2;36;24;10m█[0m[38;2;35;25;15m█[0m[38;2;14;13;9m█[0m[38;2;85;99;102m█[0m[38;2;84;95;99m█[0m[38;2;78;89;93m█[0m[38;2;88;99;103m█[0m[38;2;87;96;101m█[0m[38;2;83;92;97m█[0m[38;2;96;113;121m█[0m[38;2;93;102;107m█[0m[38;2;85;94;99m█[0m[38;2;83;92;97m█[0m[38;2;82;91;96m█[0m[38;2;78;87;92m█[0m[38;2;80;89;96m█[0m[38;2;75;85;87m█[0m[38;2;82;95;103m█[0m");
$display("[38;2;86;97;101m█[0m[38;2;99;114;121m█[0m[38;2;89;98;103m█[0m[38;2;78;87;92m█[0m[38;2;73;82;87m█[0m[38;2;77;86;91m█[0m[38;2;86;97;103m█[0m[38;2;78;89;93m█[0m[38;2;81;90;95m█[0m[38;2;80;89;94m█[0m[38;2;74;83;88m█[0m[38;2;76;85;90m█[0m[38;2;84;93;98m█[0m[38;2;80;89;94m█[0m[38;2;76;85;90m█[0m[38;2;86;99;107m█[0m[38;2;37;25;13m█[0m[38;2;11;0;0m█[0m[38;2;167;123;74m█[0m[38;2;166;126;77m█[0m[38;2;156;115;69m█[0m[38;2;158;116;74m█[0m[38;2;24;23;5m█[0m[38;2;37;15;4m█[0m[38;2;187;144;89m█[0m[38;2;182;142;83m█[0m[38;2;183;143;84m█[0m[38;2;184;142;84m█[0m[38;2;179;137;79m█[0m[38;2;182;140;82m█[0m[38;2;181;141;82m█[0m[38;2;183;143;84m█[0m[38;2;181;141;82m█[0m[38;2;178;138;79m█[0m[38;2;182;142;83m█[0m[38;2;180;140;81m█[0m[38;2;185;143;85m█[0m[38;2;188;148;89m█[0m[38;2;181;141;82m█[0m[38;2;185;143;85m█[0m[38;2;180;138;80m█[0m[38;2;180;140;81m█[0m[38;2;179;145;84m█[0m[38;2;181;141;79m█[0m[38;2;183;143;84m█[0m[38;2;186;144;86m█[0m[38;2;177;135;77m█[0m[38;2;182;140;82m█[0m[38;2;182;142;83m██[0m[38;2;209;173;125m█[0m[38;2;32;21;15m█[0m[38;2;60;46;37m█[0m[38;2;119;139;148m█[0m[38;2;110;132;145m█[0m[38;2;111;131;142m█[0m[38;2;120;145;152m█[0m[38;2;171;142;100m█[0m[38;2;185;143;85m█[0m[38;2;183;143;81m█[0m[38;2;177;141;83m█[0m[38;2;37;25;13m█[0m[38;2;33;23;14m█[0m[38;2;105;114;119m█[0m[38;2;86;99;107m█[0m[38;2;97;104;110m█[0m[38;2;97;108;114m█[0m[38;2;115;117;116m█[0m[38;2;34;24;12m█[0m[38;2;40;27;19m█[0m[38;2;176;135;79m█[0m[38;2;184;143;87m█[0m[38;2;183;143;84m█[0m[38;2;184;144;85m█[0m[38;2;183;143;84m█[0m[38;2;185;145;86m██[0m[38;2;178;138;79m█[0m[38;2;181;141;82m█[0m[38;2;182;142;83m█[0m[38;2;185;145;86m█[0m[38;2;175;135;76m█[0m[38;2;183;143;84m█[0m[38;2;180;135;78m█[0m[38;2;35;23;11m█[0m[38;2;34;23;3m█[0m[38;2;41;34;28m█[0m[38;2;102;113;117m█[0m[38;2;74;85;89m█[0m[38;2;88;99;103m█[0m[38;2;78;89;93m█[0m[38;2;83;92;97m█[0m[38;2;91;104;112m█[0m[38;2;88;96;99m█[0m[38;2;90;99;104m█[0m[38;2;83;94;98m█[0m[38;2;79;90;94m█[0m[38;2;88;99;103m█[0m[38;2;75;86;90m█[0m[38;2;89;100;104m█[0m");
$display("[38;2;92;103;107m█[0m[38;2;96;107;111m█[0m[38;2;132;149;159m█[0m[38;2;88;99;105m█[0m[38;2;89;100;102m█[0m[38;2;90;101;105m█[0m[38;2;92;102;104m█[0m[38;2;95;105;114m█[0m[38;2;88;99;103m█[0m[38;2;78;89;93m█[0m[38;2;81;92;96m█[0m[38;2;81;90;95m█[0m[38;2;85;94;99m█[0m[38;2;80;91;95m█[0m[38;2;97;108;112m█[0m[38;2;91;102;106m█[0m[38;2;31;25;11m█[0m[38;2;39;30;15m█[0m[38;2;151;119;70m█[0m[38;2;151;110;58m█[0m[38;2;183;158;118m█[0m[38;2;36;24;10m█[0m[38;2;37;28;13m█[0m[38;2;181;139;81m███[0m[38;2;182;140;82m█[0m[38;2;181;139;81m█[0m[38;2;176;134;76m█[0m[38;2;182;140;82m█[0m[38;2;185;145;86m█[0m[38;2;183;143;84m█[0m[38;2;185;145;86m█[0m[38;2;177;137;78m█[0m[38;2;175;134;78m█[0m[38;2;179;138;82m█[0m[38;2;192;152;93m█[0m[38;2;184;144;85m█[0m[38;2;183;143;84m█[0m[38;2;187;145;87m█[0m[38;2;178;136;78m█[0m[38;2;34;20;9m█[0m[38;2;81;117;149m█[0m[38;2;185;135;76m█[0m[38;2;186;144;86m█[0m[38;2;182;140;82m█[0m[38;2;185;143;85m█[0m[38;2;183;141;83m█[0m[38;2;176;134;76m█[0m[38;2;179;137;79m█[0m[38;2;187;140;84m█[0m[38;2;196;163;118m█[0m[38;2;29;25;0m█[0m[38;2;30;23;15m█[0m[38;2;39;20;5m█[0m[38;2;139;162;178m█[0m[38;2;128;145;165m█[0m[38;2;166;139;112m█[0m[38;2;182;140;82m█[0m[38;2;187;146;90m█[0m[38;2;181;139;81m█[0m[38;2;33;21;9m█[0m[38;2;32;25;6m█[0m[38;2;35;27;6m█[0m[38;2;38;21;13m█[0m[38;2;33;23;22m█[0m[38;2;39;25;14m█[0m[38;2;36;24;12m█[0m[38;2;50;36;25m█[0m[38;2;175;138;86m█[0m[38;2;181;141;82m█[0m[38;2;182;141;85m█[0m[38;2;181;141;82m█[0m[38;2;182;142;83m█[0m[38;2;186;146;87m█[0m[38;2;181;141;82m█[0m[38;2;179;139;80m█[0m[38;2;181;141;82m█[0m[38;2;178;137;81m█[0m[38;2;182;141;85m█[0m[38;2;181;141;82m██[0m[38;2;178;138;79m█[0m[38;2;180;140;81m█[0m[38;2;179;139;78m█[0m[38;2;21;2;0m█[0m[38;2;36;24;12m█[0m[38;2;37;30;22m█[0m[38;2;93;102;107m█[0m[38;2;98;107;114m█[0m[38;2;100;109;116m█[0m[38;2;84;95;99m█[0m[38;2;89;98;103m█[0m[38;2;114;131;141m█[0m[38;2;88;99;105m█[0m[38;2;95;106;110m█[0m[38;2;94;105;109m█[0m[38;2;92;103;107m█[0m[38;2;107;116;121m█[0m[38;2;89;98;103m█[0m");
$display("[38;2;99;110;114m██[0m[38;2;98;109;113m█[0m[38;2;136;153;161m█[0m[38;2;83;94;98m█[0m[38;2;97;108;112m█[0m[38;2;89;100;104m█[0m[38;2;95;106;110m█[0m[38;2;85;98;106m█[0m[38;2;93;104;110m█[0m[38;2;102;113;119m█[0m[38;2;89;100;104m█[0m[38;2;93;104;108m█[0m[38;2;89;100;104m█[0m[38;2;99;110;114m█[0m[38;2;95;106;110m█[0m[38;2;37;21;8m█[0m[38;2;39;30;15m█[0m[38;2;145;108;56m█[0m[38;2;32;22;23m█[0m[38;2;34;24;15m█[0m[38;2;185;139;87m█[0m[38;2;177;135;77m█[0m[38;2;182;143;78m█[0m[38;2;180;137;82m█[0m[38;2;180;138;80m█[0m[38;2;179;139;80m█[0m[38;2;188;146;88m█[0m[38;2;177;137;78m█[0m[38;2;185;145;86m█[0m[38;2;183;143;84m█[0m[38;2;177;135;77m██[0m[38;2;181;141;82m█[0m[38;2;186;144;86m█[0m[38;2;179;137;79m█[0m[38;2;179;139;80m█[0m[38;2;192;150;92m█[0m[38;2;180;138;80m█[0m[38;2;184;141;86m█[0m[38;2;179;138;76m█[0m[38;2;38;32;10m█[0m[38;2;90;132;154m█[0m[38;2;99;71;23m█[0m[38;2;182;137;82m█[0m[38;2;181;139;81m█[0m[38;2;183;141;83m█[0m[38;2;180;138;80m█[0m[38;2;182;140;82m█[0m[38;2;180;138;80m█[0m[38;2;183;141;83m█[0m[38;2;181;139;81m█[0m[38;2;182;140;82m█[0m[38;2;188;150;85m█[0m[38;2;182;139;70m█[0m[38;2;16;0;0m█[0m[38;2;183;140;85m█[0m[38;2;180;138;78m█[0m[38;2;179;139;80m█[0m[38;2;186;146;87m█[0m[38;2;182;140;82m█[0m[38;2;38;26;12m█[0m[38;2;29;26;7m█[0m[38;2;178;138;87m█[0m[38;2;182;140;82m█[0m[38;2;179;136;81m█[0m[38;2;183;143;82m█[0m[38;2;32;21;15m█[0m[38;2;39;22;12m█[0m[38;2;33;21;9m█[0m[38;2;37;27;17m█[0m[38;2;182;147;81m█[0m[38;2;180;140;88m█[0m[38;2;181;139;81m█[0m[38;2;183;141;83m█[0m[38;2;175;136;81m█[0m[38;2;190;140;77m█[0m[38;2;179;137;77m█[0m[38;2;185;137;71m█[0m[38;2;184;144;85m█[0m[38;2;184;147;92m█[0m[38;2;188;148;89m█[0m[38;2;180;140;81m██[0m[38;2;181;141;82m█[0m[38;2;179;139;80m█[0m[38;2;25;7;5m█[0m[38;2;34;26;15m█[0m[38;2;32;32;30m█[0m[38;2;97;108;112m█[0m[38;2;92;103;107m█[0m[38;2;88;99;103m█[0m[38;2;110;121;125m█[0m[38;2;97;108;112m█[0m[38;2;128;146;156m█[0m[38;2;93;108;115m█[0m[38;2;96;105;110m█[0m[38;2;92;101;106m█[0m[38;2;69;79;81m██[0m");
$display("[38;2;76;85;90m█[0m[38;2;75;84;89m█[0m[38;2;87;98;102m█[0m[38;2;77;87;89m█[0m[38;2;125;140;147m█[0m[38;2;117;132;139m█[0m[38;2;85;96;100m█[0m[38;2;90;101;105m█[0m[38;2;101;112;116m█[0m[38;2;88;99;105m█[0m[38;2;88;101;109m█[0m[38;2;103;114;118m█[0m[38;2;100;111;115m█[0m[38;2;99;110;116m█[0m[38;2;104;115;119m█[0m[38;2;100;111;115m█[0m[38;2;36;24;12m█[0m[38;2;35;22;13m█[0m[38;2;38;24;13m█[0m[38;2;35;28;18m█[0m[38;2;190;150;91m█[0m[38;2;184;141;86m█[0m[38;2;185;143;85m█[0m[38;2;184;142;70m█[0m[38;2;17;0;0m█[0m[38;2;90;131;151m█[0m[38;2;41;23;13m█[0m[38;2;185;139;89m█[0m[38;2;181;139;81m█[0m[38;2;182;140;82m█[0m[38;2;182;142;81m█[0m[38;2;187;145;87m█[0m[38;2;183;141;83m█[0m[38;2;180;138;80m█[0m[38;2;179;137;79m██[0m[38;2;180;140;81m█[0m[38;2;178;136;78m█[0m[38;2;183;141;83m█[0m[38;2;179;137;79m█[0m[38;2;12;2;0m█[0m[38;2;53;64;70m█[0m[38;2;81;124;156m█[0m[38;2;41;27;14m█[0m[38;2;175;135;76m█[0m[38;2;182;140;82m█[0m[38;2;181;139;81m█[0m[38;2;182;140;82m█[0m[38;2;180;138;80m█[0m[38;2;179;137;79m█[0m[38;2;182;140;82m█[0m[38;2;179;137;79m█[0m[38;2;180;138;80m█[0m[38;2;184;142;84m█[0m[38;2;181;139;81m█[0m[38;2;183;143;84m█[0m[38;2;181;141;82m█[0m[38;2;186;146;87m█[0m[38;2;179;137;79m█[0m[38;2;177;135;77m█[0m[38;2;181;139;81m█[0m[38;2;39;22;6m█[0m[38;2;31;21;11m█[0m[38;2;187;141;89m█[0m[38;2;182;142;83m█[0m[38;2;187;147;88m█[0m[38;2;183;143;84m█[0m[38;2;184;142;84m█[0m[38;2;179;137;79m█[0m[38;2;182;134;86m█[0m[38;2;32;19;0m█[0m[38;2;33;24;9m█[0m[38;2;34;22;8m█[0m[38;2;30;27;20m█[0m[38;2;176;134;84m█[0m[38;2;34;24;0m█[0m[38;2;43;28;35m█[0m[38;2;171;132;91m█[0m[38;2;137;108;76m█[0m[38;2;32;19;13m█[0m[38;2;37;26;20m█[0m[38;2;175;141;93m█[0m[38;2;184;143;87m█[0m[38;2;182;141;85m█[0m[38;2;188;148;89m█[0m[38;2;185;145;86m█[0m[38;2;182;139;88m█[0m[38;2;34;22;6m█[0m[38;2;40;24;9m█[0m[38;2;94;105;109m█[0m[38;2;95;106;110m█[0m[38;2;99;110;116m█[0m[38;2;90;103;109m█[0m[38;2;92;101;108m█[0m[38;2;104;115;117m█[0m[38;2;121;135;144m█[0m[38;2;88;99;105m█[0m[38;2;70;80;82m█[0m[38;2;71;81;83m█[0m[38;2;69;79;81m█[0m");
$display("[38;2;62;72;74m█[0m[38;2;64;74;76m█[0m[38;2;60;70;72m█[0m[38;2;62;72;74m█[0m[38;2;68;78;80m█[0m[38;2;66;75;82m█[0m[38;2;108;125;135m█[0m[38;2;62;72;74m█[0m[38;2;65;76;80m█[0m[38;2;96;107;111m█[0m[38;2;94;105;109m█[0m[38;2;109;120;126m█[0m[38;2;103;112;117m█[0m[38;2;98;109;113m█[0m[38;2;100;111;115m█[0m[38;2;97;108;112m█[0m[38;2;116;120;119m█[0m[38;2;36;24;8m█[0m[38;2;30;9;0m█[0m[38;2;181;141;82m█[0m[38;2;184;143;87m█[0m[38;2;180;139;83m█[0m[38;2;182;142;83m█[0m[38;2;187;147;88m█[0m[38;2;31;20;14m█[0m[38;2;52;66;79m█[0m[38;2;35;23;9m█[0m[38;2;181;142;85m█[0m[38;2;184;142;84m█[0m[38;2;179;137;79m█[0m[38;2;38;28;18m█[0m[38;2;84;59;28m█[0m[38;2;177;132;75m█[0m[38;2;174;144;84m█[0m[38;2;32;22;12m█[0m[38;2;190;147;69m█[0m[38;2;177;135;87m█[0m[38;2;15;0;0m█[0m[38;2;176;137;78m█[0m[38;2;184;136;90m█[0m[38;2;201;161;109m█[0m[38;2;32;22;13m█[0m[38;2;21;17;16m█[0m[38;2;39;27;15m█[0m[38;2;181;142;87m█[0m[38;2;184;142;84m██[0m[38;2;182;140;82m█[0m[38;2;181;139;81m██[0m[38;2;209;167;109m█[0m[38;2;26;5;0m█[0m[38;2;180;141;86m█[0m[38;2;180;138;80m█[0m[38;2;184;142;84m█[0m[38;2;182;142;83m█[0m[38;2;183;141;83m█[0m[38;2;187;145;87m█[0m[38;2;180;140;81m█[0m[38;2;182;140;82m█[0m[38;2;190;148;90m█[0m[38;2;188;141;87m█[0m[38;2;170;134;74m█[0m[38;2;173;134;77m█[0m[38;2;184;144;85m█[0m[38;2;180;138;80m█[0m[38;2;186;144;86m█[0m[38;2;182;140;82m█[0m[38;2;186;144;86m█[0m[38;2;177;137;78m█[0m[38;2;181;138;83m█[0m[38;2;180;139;85m█[0m[38;2;194;149;82m█[0m[38;2;29;17;5m█[0m[38;2;36;24;12m█[0m[38;2;36;20;4m█[0m[38;2;159;120;79m█[0m[38;2;156;116;67m█[0m[38;2;152;112;63m█[0m[38;2;159;119;70m█[0m[38;2;160;114;62m█[0m[38;2;34;19;12m█[0m[38;2;119;93;66m█[0m[38;2;183;142;86m█[0m[38;2;178;135;80m█[0m[38;2;186;143;88m█[0m[38;2;177;140;70m█[0m[38;2;39;27;15m█[0m[38;2;35;23;11m█[0m[38;2;112;123;127m█[0m[38;2;79;90;94m█[0m[38;2;69;79;81m█[0m[38;2;65;76;80m█[0m[38;2;66;79;85m█[0m[38;2;82;92;94m█[0m[38;2;69;78;83m█[0m[38;2;66;76;77m█[0m[38;2;59;69;71m█[0m[38;2;64;74;76m█[0m[38;2;60;70;72m█[0m");
$display("[38;2;59;69;71m█[0m[38;2;63;73;75m█[0m[38;2;74;83;88m█[0m[38;2;65;75;77m█[0m[38;2;71;81;83m█[0m[38;2;68;79;83m█[0m[38;2;58;70;70m█[0m[38;2;109;129;140m█[0m[38;2;65;75;77m█[0m[38;2;68;78;80m█[0m[38;2;66;76;78m█[0m[38;2;62;72;74m█[0m[38;2;68;78;80m█[0m[38;2;71;82;84m█[0m[38;2;98;109;113m█[0m[38;2;96;107;111m█[0m[38;2;35;23;11m█[0m[38;2;42;21;18m█[0m[38;2;186;146;85m█[0m[38;2;184;143;87m█[0m[38;2;186;146;87m█[0m[38;2;184;144;85m█[0m[38;2;182;140;82m█[0m[38;2;192;140;90m█[0m[38;2;186;138;89m█[0m[38;2;185;138;82m█[0m[38;2;184;145;90m█[0m[38;2;184;136;74m█[0m[38;2;206;174;136m█[0m[38;2;39;21;19m█[0m[38;2;207;174;133m█[0m[38;2;185;144;90m█[0m[38;2;178;136;78m█[0m[38;2;178;139;70m█[0m[38;2;20;17;10m█[0m[38;2;12;0;0m█[0m[38;2;182;132;83m█[0m[38;2;30;24;2m█[0m[38;2;32;21;17m█[0m[38;2;181;139;81m█[0m[38;2;184;142;84m█[0m[38;2;178;139;74m█[0m[38;2;176;133;78m█[0m[38;2;186;141;82m█[0m[38;2;180;138;80m█[0m[38;2;184;142;84m█[0m[38;2;185;143;85m█[0m[38;2;184;142;84m█[0m[38;2;189;149;90m█[0m[38;2;181;139;81m█[0m[38;2;37;25;11m█[0m[38;2;106;150;189m█[0m[38;2;102;139;158m█[0m[38;2;202;169;134m█[0m[38;2;180;138;80m█[0m[38;2;181;139;81m█[0m[38;2;184;142;84m█[0m[38;2;185;143;85m█[0m[38;2;177;137;78m█[0m[38;2;179;137;79m█[0m[38;2;182;140;82m█[0m[38;2;183;143;84m█[0m[38;2;188;150;88m█[0m[38;2;29;29;19m█[0m[38;2;174;137;84m█[0m[38;2;191;150;98m█[0m[38;2;183;143;84m█[0m[38;2;181;141;82m█[0m[38;2;185;145;86m█[0m[38;2;181;141;82m█[0m[38;2;179;137;79m█[0m[38;2;179;139;80m█[0m[38;2;177;137;78m█[0m[38;2;183;147;87m█[0m[38;2;172;138;67m█[0m[38;2;33;19;8m█[0m[38;2;36;22;11m█[0m[38;2;13;0;0m█[0m[38;2;159;119;70m█[0m[38;2;153;113;64m█[0m[38;2;147;112;56m█[0m[38;2;38;26;10m█[0m[38;2;40;25;2m█[0m[38;2;155;114;68m█[0m[38;2;157;116;70m█[0m[38;2;155;114;68m█[0m[38;2;155;116;75m█[0m[38;2;39;25;14m█[0m[38;2;36;22;11m█[0m[38;2;64;75;79m█[0m[38;2;67;78;82m█[0m[38;2;72;82;84m█[0m[38;2;62;73;75m█[0m[38;2;54;67;73m█[0m[38;2;115;130;135m█[0m[38;2;63;73;75m█[0m[38;2;70;80;82m█[0m[38;2;62;72;74m█[0m[38;2;63;71;74m█[0m[38;2;69;77;80m█[0m");
$display("[38;2;63;71;74m█[0m[38;2;60;68;71m██[0m[38;2;97;110;116m█[0m[38;2;60;65;71m█[0m[38;2;63;71;74m█[0m[38;2;58;68;70m█[0m[38;2;59;69;71m█[0m[38;2;98;108;117m█[0m[38;2;65;73;76m█[0m[38;2;68;76;79m█[0m[38;2;66;76;78m█[0m[38;2;61;71;73m██[0m[38;2;60;73;79m█[0m[38;2;41;27;14m█[0m[38;2;30;23;17m█[0m[38;2;183;143;84m█[0m[38;2;188;148;89m█[0m[38;2;177;137;78m█[0m[38;2;185;143;85m█[0m[38;2;181;139;81m█[0m[38;2;180;140;81m█[0m[38;2;180;141;82m█[0m[38;2;183;143;84m█[0m[38;2;181;141;82m█[0m[38;2;179;139;80m█[0m[38;2;181;141;82m█[0m[38;2;186;144;86m█[0m[38;2;181;139;81m█[0m[38;2;182;140;82m█[0m[38;2;189;147;89m█[0m[38;2;183;141;83m█[0m[38;2;186;144;86m█[0m[38;2;187;147;88m█[0m[38;2;187;145;87m█[0m[38;2;183;143;84m█[0m[38;2;189;147;89m█[0m[38;2;185;143;85m█[0m[38;2;180;138;80m█[0m[38;2;183;141;83m█[0m[38;2;176;134;76m█[0m[38;2;181;139;81m█[0m[38;2;179;137;79m█[0m[38;2;181;139;81m█[0m[38;2;174;132;74m█[0m[38;2;184;142;84m█[0m[38;2;177;135;77m█[0m[38;2;185;143;85m█[0m[38;2;178;136;78m█[0m[38;2;34;21;5m█[0m[38;2;137;154;162m█[0m[38;2;54;72;82m█[0m[38;2;40;30;20m█[0m[38;2;186;142;81m█[0m[38;2;182;140;82m█[0m[38;2;177;136;80m█[0m[38;2;189;148;92m█[0m[38;2;184;144;85m█[0m[38;2;182;140;82m█[0m[38;2;194;152;94m█[0m[38;2;188;146;88m█[0m[38;2;182;142;83m█[0m[38;2;204;154;101m█[0m[38;2;37;20;4m█[0m[38;2;178;129;70m█[0m[38;2;174;133;79m█[0m[38;2;185;143;85m█[0m[38;2;181;139;81m█[0m[38;2;183;141;83m███[0m[38;2;183;143;84m█[0m[38;2;184;142;84m█[0m[38;2;181;139;81m█[0m[38;2;191;149;91m█[0m[38;2;203;161;103m█[0m[38;2;40;26;13m█[0m[38;2;36;25;3m█[0m[38;2;166;120;61m█[0m[38;2;158;107;64m█[0m[38;2;33;24;9m█[0m[38;2;20;0;0m█[0m[38;2;158;118;69m█[0m[38;2;158;118;67m█[0m[38;2;153;113;64m█[0m[38;2;28;6;0m█[0m[38;2;36;22;11m█[0m[38;2;24;11;5m█[0m[38;2;61;71;73m█[0m[38;2;64;74;76m█[0m[38;2;58;68;70m█[0m[38;2;64;72;75m█[0m[38;2;68;76;79m█[0m[38;2;59;67;69m█[0m[38;2;93;109;122m█[0m[38;2;56;67;69m█[0m[38;2;51;59;62m█[0m[38;2;57;65;67m██[0m");
$display("[38;2;59;67;70m█[0m[38;2;61;69;72m█[0m[38;2;63;71;74m█[0m[38;2;60;70;72m█[0m[38;2;89;103;112m█[0m[38;2;65;75;76m█[0m[38;2;61;69;72m█[0m[38;2;66;74;77m█[0m[38;2;58;66;69m█[0m[38;2;73;81;84m█[0m[38;2;65;73;76m███[0m[38;2;64;72;75m█[0m[38;2;72;71;66m█[0m[38;2;34;22;10m█[0m[38;2;178;158;123m█[0m[38;2;186;146;87m█[0m[38;2;178;138;79m█[0m[38;2;181;141;82m█[0m[38;2;182;140;82m█[0m[38;2;180;138;80m█[0m[38;2;186;146;87m█[0m[38;2;179;137;79m█[0m[38;2;180;138;80m█[0m[38;2;184;141;86m█[0m[38;2;183;140;85m█[0m[38;2;184;142;84m█[0m[38;2;179;139;80m█[0m[38;2;182;142;83m█[0m[38;2;185;143;85m█[0m[38;2;183;143;84m██[0m[38;2;175;135;76m█[0m[38;2;182;140;82m█[0m[38;2;185;143;85m█[0m[38;2;186;146;87m█[0m[38;2;179;137;79m█[0m[38;2;183;141;83m█[0m[38;2;182;141;87m█[0m[38;2;178;135;80m█[0m[38;2;186;144;86m█[0m[38;2;188;146;88m█[0m[38;2;185;143;85m█[0m[38;2;174;132;74m█[0m[38;2;188;147;91m█[0m[38;2;180;138;80m█[0m[38;2;189;147;89m█[0m[38;2;183;141;83m█[0m[38;2;181;139;81m█[0m[38;2;182;134;86m█[0m[38;2;20;0;0m█[0m[38;2;200;165;125m█[0m[38;2;181;139;81m█[0m[38;2;183;141;83m█[0m[38;2;183;143;84m█[0m[38;2;184;142;84m█[0m[38;2;183;141;83m█[0m[38;2;178;138;79m█[0m[38;2;182;142;83m█[0m[38;2;180;140;81m█[0m[38;2;185;143;85m█[0m[38;2;185;142;87m█[0m[38;2;178;136;78m█[0m[38;2;36;18;4m█[0m[38;2;32;24;11m█[0m[38;2;179;143;83m█[0m[38;2;182;142;83m█[0m[38;2;178;138;79m█[0m[38;2;189;147;89m█[0m[38;2;59;37;16m█[0m[38;2;175;138;83m█[0m[38;2;183;141;83m█[0m[38;2;178;138;79m█[0m[38;2;184;144;85m█[0m[38;2;185;145;86m█[0m[38;2;186;146;87m█[0m[38;2;179;139;78m█[0m[38;2;33;23;13m█[0m[38;2;35;22;13m█[0m[38;2;32;24;13m█[0m[38;2;19;0;0m█[0m[38;2;144;103;57m█[0m[38;2;158;118;69m█[0m[38;2;153;113;62m█[0m[38;2;148;118;94m█[0m[38;2;36;24;12m█[0m[38;2;33;19;6m█[0m[38;2;63;73;75m█[0m[38;2;66;76;78m██[0m[38;2;60;70;72m█[0m[38;2;52;60;62m█[0m[38;2;53;61;63m█[0m[38;2;50;58;60m█[0m[38;2;56;66;67m█[0m[38;2;82;97;104m█[0m[38;2;50;58;61m█[0m[38;2;46;54;56m█[0m[38;2;44;52;54m█[0m");
$display("[38;2;46;54;56m█[0m[38;2;44;52;54m█[0m[38;2;50;58;60m█[0m[38;2;53;61;64m█[0m[38;2;65;73;76m█[0m[38;2;99;116;126m█[0m[38;2;60;70;72m█[0m[38;2;59;67;70m█[0m[38;2;52;60;62m█[0m[38;2;50;58;60m█[0m[38;2;48;56;58m█[0m[38;2;53;61;64m█[0m[38;2;65;73;76m█[0m[38;2;55;63;66m█[0m[38;2;35;22;14m█[0m[38;2;36;22;11m█[0m[38;2;179;142;89m█[0m[38;2;181;141;82m█[0m[38;2;183;143;84m█[0m[38;2;182;142;83m█[0m[38;2;183;149;112m█[0m[38;2;35;27;4m█[0m[38;2;40;21;7m█[0m[38;2;36;18;8m█[0m[38;2;42;23;17m█[0m[38;2;33;21;5m█[0m[38;2;31;19;0m█[0m[38;2;35;23;11m█[0m[38;2;26;18;5m█[0m[38;2;189;146;91m█[0m[38;2;181;139;81m█[0m[38;2;181;141;82m█[0m[38;2;178;138;79m█[0m[38;2;178;136;78m█[0m[38;2;184;144;85m█[0m[38;2;183;143;84m█[0m[38;2;181;139;81m█[0m[38;2;182;142;83m█[0m[38;2;185;145;86m█[0m[38;2;35;25;16m█[0m[38;2;37;25;11m█[0m[38;2;30;18;6m█[0m[38;2;39;21;9m█[0m[38;2;43;25;11m█[0m[38;2;39;20;6m█[0m[38;2;38;28;16m█[0m[38;2;31;22;7m█[0m[38;2;38;28;16m█[0m[38;2;30;4;0m█[0m[38;2;185;143;83m█[0m[38;2;183;141;83m█[0m[38;2;185;143;85m█[0m[38;2;181;139;81m█[0m[38;2;177;135;77m█[0m[38;2;191;149;91m█[0m[38;2;182;142;83m█[0m[38;2;186;146;87m█[0m[38;2;178;138;79m█[0m[38;2;194;148;88m█[0m[38;2;144;142;143m█[0m[38;2;184;138;78m█[0m[38;2;186;144;86m█[0m[38;2;180;140;81m█[0m[38;2;188;148;89m█[0m[38;2;195;158;103m█[0m[38;2;34;22;6m█[0m[38;2;208;176;115m█[0m[38;2;184;141;86m█[0m[38;2;183;140;85m█[0m[38;2;181;142;77m█[0m[38;2;28;19;4m█[0m[38;2;73;128;169m█[0m[38;2;176;145;80m█[0m[38;2;182;142;83m█[0m[38;2;187;147;88m█[0m[38;2;180;140;81m█[0m[38;2;178;138;79m█[0m[38;2;182;140;82m█[0m[38;2;182;135;83m█[0m[38;2;42;24;10m█[0m[38;2;33;20;11m█[0m[38;2;155;115;66m█[0m[38;2;155;114;68m█[0m[38;2;156;119;64m█[0m[38;2;45;33;19m█[0m[38;2;35;23;11m█[0m[38;2;34;24;14m█[0m[38;2;66;74;77m█[0m[38;2;58;66;69m█[0m[38;2;59;67;70m█[0m[38;2;54;62;65m█[0m[38;2;72;83;87m█[0m[38;2;47;55;57m█[0m[38;2;51;59;61m█[0m[38;2;49;57;59m█[0m[38;2;50;58;60m█[0m[38;2;53;61;63m█[0m[38;2;44;52;54m█[0m[38;2;49;57;59m██[0m");
$display("[38;2;45;53;55m█[0m[38;2;48;56;58m█[0m[38;2;51;59;61m█[0m[38;2;49;57;59m█[0m[38;2;47;55;57m█[0m[38;2;54;63;62m█[0m[38;2;95;109;118m█[0m[38;2;46;56;57m█[0m[38;2;47;55;57m█[0m[38;2;49;57;59m█[0m[38;2;56;64;66m█[0m[38;2;48;56;58m██[0m[38;2;55;65;67m█[0m[38;2;35;23;11m█[0m[38;2;39;27;15m█[0m[38;2;170;125;70m█[0m[38;2;181;141;82m█[0m[38;2;177;137;78m█[0m[38;2;179;137;79m█[0m[38;2;176;139;86m█[0m[38;2;184;141;86m█[0m[38;2;180;138;78m█[0m[38;2;185;140;83m█[0m[38;2;181;139;81m█[0m[38;2;180;141;82m█[0m[38;2;191;149;101m█[0m[38;2;187;148;89m█[0m[38;2;180;138;80m█[0m[38;2;181;139;81m█[0m[38;2;178;133;74m█[0m[38;2;181;143;94m█[0m[38;2;195;146;79m█[0m[38;2;188;137;80m█[0m[38;2;185;138;82m█[0m[38;2;182;140;90m█[0m[38;2;178;138;79m█[0m[38;2;182;140;82m█[0m[38;2;184;142;84m█[0m[38;2;176;135;79m█[0m[38;2;183;138;79m█[0m[38;2;184;142;82m█[0m[38;2;186;143;75m█[0m[38;2;187;144;93m█[0m[38;2;177;139;77m█[0m[38;2;179;145;84m█[0m[38;2;176;141;87m█[0m[38;2;188;149;94m█[0m[38;2;187;145;85m█[0m[38;2;185;141;92m█[0m[38;2;188;148;89m█[0m[38;2;187;147;88m█[0m[38;2;183;143;84m█[0m[38;2;182;140;82m█[0m[38;2;186;144;86m█[0m[38;2;182;142;83m█[0m[38;2;181;139;81m█[0m[38;2;180;138;80m█[0m[38;2;178;131;85m█[0m[38;2;35;18;8m█[0m[38;2;137;145;106m█[0m[38;2;185;143;85m█[0m[38;2;177;135;77m█[0m[38;2;180;138;80m█[0m[38;2;177;140;85m█[0m[38;2;35;23;11m█[0m[38;2;25;22;17m█[0m[38;2;182;140;82m█[0m[38;2;181;139;81m█[0m[38;2;177;138;81m█[0m[38;2;35;22;13m█[0m[38;2;96;131;159m█[0m[38;2;44;23;28m█[0m[38;2;184;142;84m█[0m[38;2;186;144;86m█[0m[38;2;181;141;82m█[0m[38;2;176;136;77m█[0m[38;2;185;143;85m█[0m[38;2;176;135;81m█[0m[38;2;186;141;82m█[0m[38;2;31;22;17m█[0m[38;2;36;22;13m█[0m[38;2;37;23;12m█[0m[38;2;35;23;11m█[0m[38;2;40;27;18m█[0m[38;2;60;70;72m█[0m[38;2;58;66;69m█[0m[38;2;53;61;64m█[0m[38;2;59;67;70m█[0m[38;2;52;60;62m█[0m[38;2;57;65;67m█[0m[38;2;53;61;63m█[0m[38;2;99;112;118m█[0m[38;2;57;65;68m█[0m[38;2;52;60;62m█[0m[38;2;49;57;59m█[0m[38;2;51;59;61m█[0m[38;2;48;56;58m█[0m[38;2;50;58;60m██[0m");
$display("[38;2;47;55;57m█[0m[38;2;48;56;58m█[0m[38;2;54;59;62m█[0m[38;2;47;55;57m█[0m[38;2;48;56;59m█[0m[38;2;50;58;60m█[0m[38;2;47;57;58m█[0m[38;2;63;74;76m█[0m[38;2;41;51;52m█[0m[38;2;47;55;57m█[0m[38;2;48;56;58m█[0m[38;2;55;63;65m█[0m[38;2;48;56;58m█[0m[38;2;36;20;7m██[0m[38;2;187;144;93m█[0m[38;2;183;143;84m█[0m[38;2;184;144;83m█[0m[38;2;179;140;85m█[0m[38;2;190;150;91m█[0m[38;2;73;51;10m█[0m[38;2;33;24;15m█[0m[38;2;36;21;16m█[0m[38;2;34;22;10m█[0m[38;2;38;26;14m█[0m[38;2;35;23;11m█[0m[38;2;39;25;16m█[0m[38;2;33;23;14m█[0m[38;2;237;229;210m█[0m[38;2;221;210;190m█[0m[38;2;224;214;187m█[0m[38;2;227;215;191m█[0m[38;2;226;214;190m█[0m[38;2;228;216;192m█[0m[38;2;224;212;188m██[0m[38;2;220;213;187m█[0m[38;2;212;207;177m█[0m[38;2;238;218;193m█[0m[38;2;204;167;123m█[0m[38;2;35;18;2m█[0m[38;2;33;19;6m█[0m[38;2;39;22;14m█[0m[38;2;38;24;11m█[0m[38;2;41;29;17m█[0m[38;2;32;24;13m█[0m[38;2;30;22;11m█[0m[38;2;40;21;7m█[0m[38;2;51;17;0m█[0m[38;2;184;141;86m█[0m[38;2;178;138;79m█[0m[38;2;182;142;83m█[0m[38;2;184;142;84m█[0m[38;2;182;140;82m█[0m[38;2;185;152;99m█[0m[38;2;171;127;64m█[0m[38;2;175;129;70m█[0m[38;2;185;135;72m█[0m[38;2;40;27;21m█[0m[38;2;123;152;170m█[0m[38;2;93;139;173m█[0m[38;2;38;27;21m█[0m[38;2;182;140;82m█[0m[38;2;188;146;88m█[0m[38;2;179;142;89m█[0m[38;2;35;23;11m█[0m[38;2;35;30;36m█[0m[38;2;184;142;84m██[0m[38;2;176;145;81m█[0m[38;2;37;23;14m█[0m[38;2;84;128;163m█[0m[38;2;29;26;11m█[0m[38;2;179;137;79m█[0m[38;2;178;136;78m█[0m[38;2;177;137;78m█[0m[38;2;183;143;84m█[0m[38;2;179;137;79m█[0m[38;2;183;143;84m█[0m[38;2;181;141;82m█[0m[38;2;201;165;107m█[0m[38;2;44;32;20m█[0m[38;2;33;21;9m█[0m[38;2;59;68;73m█[0m[38;2;62;70;73m█[0m[38;2;57;65;68m█[0m[38;2;53;61;63m█[0m[38;2;48;56;58m█[0m[38;2;46;54;56m█[0m[38;2;48;56;58m███[0m[38;2;52;60;62m█[0m[38;2;74;90;103m█[0m[38;2;54;62;65m█[0m[38;2;49;57;59m█[0m[38;2;47;55;57m█[0m[38;2;42;50;52m█[0m[38;2;45;53;55m█[0m[38;2;44;52;54m█[0m");
$display("[38;2;54;53;48m██[0m[38;2;51;50;46m█[0m[38;2;48;47;42m█[0m[38;2;48;48;46m█[0m[38;2;50;51;46m█[0m[38;2;56;53;48m█[0m[38;2;51;48;43m█[0m[38;2;53;52;47m█[0m[38;2;49;49;41m█[0m[38;2;50;50;42m█[0m[38;2;52;49;42m█[0m[38;2;20;15;9m█[0m[38;2;33;24;17m█[0m[38;2;162;128;65m█[0m[38;2;228;209;177m█[0m[38;2;227;212;183m█[0m[38;2;227;215;191m█[0m[38;2;229;221;200m█[0m[38;2;228;216;192m█[0m[38;2;220;214;192m█[0m[38;2;227;217;192m█[0m[38;2;223;211;195m█[0m[38;2;228;217;189m█[0m[38;2;231;214;184m█[0m[38;2;229;214;185m█[0m[38;2;222;214;193m█[0m[38;2;223;213;188m█[0m[38;2;255;252;231m█[0m[38;2;34;22;6m█[0m[38;2;34;24;14m█[0m[38;2;34;24;12m██[0m[38;2;38;24;13m█[0m[38;2;36;27;18m█[0m[38;2;225;213;189m█[0m[38;2;231;219;195m█[0m[38;2;225;213;189m█[0m[38;2;230;218;194m█[0m[38;2;222;214;191m█[0m[38;2;226;211;182m█[0m[38;2;229;213;190m█[0m[38;2;248;232;199m█[0m[38;2;200;150;87m█[0m[38;2;186;145;93m█[0m[38;2;187;155;96m█[0m[38;2;169;137;76m█[0m[38;2;177;135;75m█[0m[38;2;154;117;62m█[0m[38;2;220;213;185m█[0m[38;2;224;216;193m█[0m[38;2;230;213;195m█[0m[38;2;222;209;192m█[0m[38;2;221;209;183m█[0m[38;2;225;214;192m█[0m[38;2;221;209;185m█[0m[38;2;228;216;192m█[0m[38;2;229;217;193m█[0m[38;2;41;28;19m█[0m[38;2;0;2;9m█[0m[38;2;139;174;202m█[0m[38;2;38;28;16m█[0m[38;2;234;194;135m█[0m[38;2;179;139;80m█[0m[38;2;236;185;119m█[0m[38;2;39;22;4m█[0m[38;2;91;70;41m█[0m[38;2;184;142;84m█[0m[38;2;181;139;81m█[0m[38;2;183;142;78m█[0m[38;2;178;138;79m█[0m[38;2;37;24;16m█[0m[38;2;210;179;150m█[0m[38;2;182;140;82m█[0m[38;2;180;138;80m█[0m[38;2;177;137;78m█[0m[38;2;191;151;92m█[0m[38;2;180;138;80m█[0m[38;2;177;138;81m█[0m[38;2;181;142;85m█[0m[38;2;189;137;79m█[0m[38;2;41;28;20m█[0m[38;2;33;20;11m█[0m[38;2;36;26;16m█[0m[38;2;39;26;10m█[0m[38;2;62;61;56m█[0m[38;2;52;49;44m█[0m[38;2;54;51;46m█[0m[38;2;51;48;43m█[0m[38;2;57;54;49m█[0m[38;2;56;53;48m█[0m[38;2;50;47;42m█[0m[38;2;54;53;48m█[0m[38;2;54;51;44m█[0m[38;2;107;129;142m█[0m[38;2;49;48;43m█[0m[38;2;51;50;45m█[0m[38;2;52;51;46m███[0m");
$display("[38;2;49;49;47m█[0m[38;2;51;51;49m█[0m[38;2;51;50;45m█[0m[38;2;49;48;43m█[0m[38;2;53;52;47m█[0m[38;2;56;55;50m█[0m[38;2;46;50;49m█[0m[38;2;52;53;47m█[0m[38;2;53;50;45m██[0m[38;2;51;48;43m█[0m[38;2;50;47;42m█[0m[38;2;37;22;17m█[0m[38;2;8;0;0m█[0m[38;2;226;214;190m██[0m[38;2;224;213;191m█[0m[38;2;223;205;195m█[0m[38;2;228;213;172m█[0m[38;2;224;212;188m█[0m[38;2;226;214;190m█[0m[38;2;225;213;189m█[0m[38;2;224;214;189m█[0m[38;2;229;217;193m█[0m[38;2;226;214;190m█[0m[38;2;225;213;189m█[0m[38;2;227;215;191m█[0m[38;2;226;214;190m█[0m[38;2;9;0;0m█[0m[38;2;35;23;11m█[0m[38;2;34;22;10m██[0m[38;2;36;24;12m█[0m[38;2;36;24;10m█[0m[38;2;27;16;10m█[0m[38;2;220;210;185m█[0m[38;2;225;213;189m██[0m[38;2;229;217;193m█[0m[38;2;223;211;187m█[0m[38;2;225;213;189m█[0m[38;2;227;215;191m█[0m[38;2;225;213;189m██[0m[38;2;227;215;191m█[0m[38;2;226;214;190m██[0m[38;2;225;213;189m█[0m[38;2;225;213;187m█[0m[38;2;225;213;191m█[0m[38;2;222;210;186m█[0m[38;2;228;216;192m█[0m[38;2;226;214;190m█[0m[38;2;223;211;187m██[0m[38;2;224;212;188m██[0m[38;2;223;211;187m█[0m[38;2;224;212;188m█[0m[38;2;255;252;233m█[0m[38;2;255;255;236m█[0m[38;2;225;213;189m█[0m[38;2;225;215;188m█[0m[38;2;226;216;189m█[0m[38;2;35;22;13m█[0m[38;2;37;25;13m█[0m[38;2;180;147;76m█[0m[38;2;187;147;88m█[0m[38;2;184;142;84m█[0m[38;2;183;141;83m█[0m[38;2;188;146;88m█[0m[38;2;179;137;79m█[0m[38;2;183;143;84m█[0m[38;2;179;139;80m█[0m[38;2;183;143;84m█[0m[38;2;185;143;85m██[0m[38;2;183;143;84m██[0m[38;2;187;147;88m█[0m[38;2;178;138;79m█[0m[38;2;190;144;95m█[0m[38;2;38;21;14m█[0m[38;2;220;212;189m█[0m[38;2;163;157;145m█[0m[38;2;37;24;15m█[0m[38;2;38;24;11m█[0m[38;2;33;21;9m█[0m[38;2;48;45;40m█[0m[38;2;53;50;43m█[0m[38;2;46;46;38m█[0m[38;2;48;47;42m█[0m[38;2;54;53;48m█[0m[38;2;47;46;41m█[0m[38;2;51;51;43m█[0m[38;2;83;102;116m█[0m[38;2;53;48;42m█[0m[38;2;56;53;48m█[0m[38;2;47;46;41m█[0m[38;2;49;48;43m█[0m");
$display("[38;2;43;44;38m█[0m[38;2;91;101;111m█[0m[38;2;47;48;42m█[0m[38;2;49;48;43m█[0m[38;2;46;45;40m█[0m[38;2;48;47;42m█[0m[38;2;49;48;43m█[0m[38;2;46;45;41m█[0m[38;2;44;43;38m█[0m[38;2;57;54;49m█[0m[38;2;53;50;45m█[0m[38;2;45;38;28m█[0m[38;2;35;23;11m█[0m[38;2;219;213;189m█[0m[38;2;224;212;188m██[0m[38;2;255;250;233m█[0m[38;2;114;151;178m█[0m[38;2;219;214;194m█[0m[38;2;224;213;191m█[0m[38;2;227;216;194m█[0m[38;2;226;215;193m█[0m[38;2;225;213;189m█[0m[38;2;226;214;190m█[0m[38;2;224;212;188m█[0m[38;2;226;214;190m█[0m[38;2;225;213;189m█[0m[38;2;223;211;187m█[0m[38;2;226;214;190m█[0m[38;2;221;209;185m█[0m[38;2;221;216;196m█[0m[38;2;34;22;8m█[0m[38;2;249;239;227m█[0m[38;2;228;218;193m█[0m[38;2;226;214;190m█[0m[38;2;227;215;191m█[0m[38;2;225;213;189m█[0m[38;2;226;214;190m█[0m[38;2;224;212;186m█[0m[38;2;228;216;192m█[0m[38;2;226;214;190m█[0m[38;2;228;216;192m█[0m[38;2;225;213;189m██[0m[38;2;228;216;192m█[0m[38;2;226;214;190m██[0m[38;2;225;213;191m█[0m[38;2;226;214;190m█[0m[38;2;229;217;193m█[0m[38;2;226;214;192m█[0m[38;2;215;206;189m█[0m[38;2;38;31;25m█[0m[38;2;229;217;191m█[0m[38;2;225;210;187m█[0m[38;2;226;214;190m█[0m[38;2;225;213;189m█[0m[38;2;222;210;186m█[0m[38;2;223;211;187m█[0m[38;2;224;212;188m█[0m[38;2;228;216;192m█[0m[38;2;227;215;191m█[0m[38;2;231;216;197m█[0m[38;2;8;0;0m█[0m[38;2;38;27;9m█[0m[38;2;173;140;105m█[0m[38;2;183;143;84m█[0m[38;2;183;141;83m█[0m[38;2;182;140;82m█[0m[38;2;179;139;80m█[0m[38;2;184;142;84m█[0m[38;2;182;140;82m█[0m[38;2;181;141;82m██[0m[38;2;182;142;83m█[0m[38;2;179;140;85m█[0m[38;2;185;139;80m█[0m[38;2;176;135;79m█[0m[38;2;176;136;77m█[0m[38;2;180;140;81m██[0m[38;2;179;138;82m█[0m[38;2;163;135;95m█[0m[38;2;221;211;186m█[0m[38;2;227;215;191m█[0m[38;2;223;211;187m█[0m[38;2;227;217;192m█[0m[38;2;8;0;0m█[0m[38;2;33;21;9m█[0m[38;2;35;23;11m█[0m[38;2;39;30;21m█[0m[38;2;46;47;41m█[0m[38;2;46;47;42m█[0m[38;2;43;44;39m█[0m[38;2;44;43;39m█[0m[38;2;44;45;40m█[0m[38;2;41;42;37m█[0m[38;2;45;46;41m█[0m[38;2;48;49;44m█[0m[38;2;46;47;42m█[0m");
$display("[38;2;56;55;50m█[0m[38;2;59;58;53m█[0m[38;2;79;96;106m█[0m[38;2;52;51;46m█[0m[38;2;51;50;45m██[0m[38;2;55;54;49m█[0m[38;2;43;42;38m█[0m[38;2;48;47;43m█[0m[38;2;53;52;47m█[0m[38;2;44;43;38m█[0m[38;2;59;54;48m█[0m[38;2;34;21;13m█[0m[38;2;251;243;224m█[0m[38;2;218;208;183m█[0m[38;2;222;210;186m█[0m[38;2;35;25;15m█[0m[38;2;82;125;157m█[0m[38;2;40;58;70m█[0m[38;2;218;207;185m█[0m[38;2;228;216;192m█[0m[38;2;224;212;188m█[0m[38;2;223;211;187m█[0m[38;2;227;215;191m█[0m[38;2;225;213;189m█[0m[38;2;224;214;189m█[0m[38;2;225;215;190m█[0m[38;2;226;214;190m█[0m[38;2;225;210;187m█[0m[38;2;223;213;188m█[0m[38;2;111;101;91m█[0m[38;2;34;24;12m█[0m[38;2;38;28;19m█[0m[38;2;214;206;187m█[0m[38;2;231;219;195m█[0m[38;2;221;209;187m█[0m[38;2;229;219;194m█[0m[38;2;227;215;191m█[0m[38;2;226;214;190m█[0m[38;2;224;212;188m█[0m[38;2;225;213;189m█[0m[38;2;224;212;188m█[0m[38;2;223;213;188m█[0m[38;2;226;216;191m█[0m[38;2;229;217;193m█[0m[38;2;223;211;187m█[0m[38;2;224;212;188m█[0m[38;2;227;215;191m█[0m[38;2;226;216;191m█[0m[38;2;223;213;188m█[0m[38;2;228;214;188m█[0m[38;2;32;18;9m█[0m[38;2;99;142;177m█[0m[38;2;29;20;5m█[0m[38;2;220;208;186m█[0m[38;2;226;214;190m█[0m[38;2;227;215;191m██[0m[38;2;221;209;185m█[0m[38;2;223;211;187m█[0m[38;2;225;213;189m█[0m[38;2;226;214;188m█[0m[38;2;28;18;8m█[0m[38;2;35;21;10m█[0m[38;2;68;45;4m█[0m[38;2;179;140;81m█[0m[38;2;179;137;79m█[0m[38;2;179;139;80m██[0m[38;2;184;142;84m█[0m[38;2;187;147;88m█[0m[38;2;177;137;78m█[0m[38;2;183;143;84m█[0m[38;2;187;145;87m█[0m[38;2;179;137;79m█[0m[38;2;184;144;93m█[0m[38;2;36;19;25m█[0m[38;2;185;152;101m█[0m[38;2;182;142;83m█[0m[38;2;184;144;85m█[0m[38;2;181;141;82m█[0m[38;2;178;138;79m█[0m[38;2;177;137;78m█[0m[38;2;235;221;195m█[0m[38;2;228;216;192m█[0m[38;2;225;213;189m█[0m[38;2;220;210;185m█[0m[38;2;226;214;190m█[0m[38;2;223;211;187m█[0m[38;2;224;213;193m█[0m[38;2;37;25;11m█[0m[38;2;31;19;7m█[0m[38;2;54;53;48m█[0m[38;2;54;51;44m█[0m[38;2;51;50;45m█[0m[38;2;53;50;45m█[0m[38;2;48;45;40m█[0m[38;2;51;48;43m█[0m[38;2;50;47;42m█[0m[38;2;53;50;45m█[0m");
$display("[38;2;52;51;46m█[0m[38;2;56;55;50m█[0m[38;2;59;56;51m█[0m[38;2;89;106;116m█[0m[38;2;51;51;43m█[0m[38;2;51;50;45m█[0m[38;2;49;48;44m█[0m[38;2;53;52;48m█[0m[38;2;50;49;45m█[0m[38;2;47;46;42m█[0m[38;2;54;53;49m█[0m[38;2;53;52;47m█[0m[38;2;39;27;15m█[0m[38;2;32;19;10m█[0m[38;2;218;211;185m█[0m[38;2;227;215;193m█[0m[38;2;31;21;12m█[0m[38;2;73;81;100m█[0m[38;2;34;22;6m█[0m[38;2;242;235;216m█[0m[38;2;225;215;190m█[0m[38;2;224;214;189m█[0m[38;2;226;214;190m█[0m[38;2;224;214;189m█[0m[38;2;222;212;187m█[0m[38;2;225;215;190m██[0m[38;2;37;27;15m█[0m[38;2;40;28;16m█[0m[38;2;34;24;12m█[0m[38;2;23;11;0m█[0m[38;2;154;105;98m█[0m[38;2;45;32;23m█[0m[38;2;37;31;17m█[0m[38;2;30;18;6m█[0m[38;2;39;25;12m█[0m[38;2;37;25;11m█[0m[38;2;29;20;11m█[0m[38;2;255;255;236m█[0m[38;2;224;212;188m█[0m[38;2;225;213;189m█[0m[38;2;223;213;188m█[0m[38;2;228;216;192m█[0m[38;2;223;211;187m█[0m[38;2;224;212;188m█[0m[38;2;221;209;185m█[0m[38;2;225;213;189m██[0m[38;2;229;217;193m█[0m[38;2;222;210;186m█[0m[38;2;224;212;188m█[0m[38;2;25;16;7m█[0m[38;2;37;24;8m█[0m[38;2;44;32;20m█[0m[38;2;225;213;187m█[0m[38;2;227;215;191m██[0m[38;2;226;214;190m█[0m[38;2;223;211;187m█[0m[38;2;222;210;188m█[0m[38;2;220;210;185m█[0m[38;2;35;23;11m█[0m[38;2;31;24;16m█[0m[38;2;192;145;93m█[0m[38;2;187;147;88m█[0m[38;2;179;139;80m█[0m[38;2;182;142;83m█[0m[38;2;183;141;83m█[0m[38;2;184;142;84m██[0m[38;2;179;137;79m█[0m[38;2;183;141;83m█[0m[38;2;178;138;79m█[0m[38;2;180;140;81m█[0m[38;2;187;147;88m█[0m[38;2;202;165;113m█[0m[38;2;34;26;5m█[0m[38;2;88;128;153m█[0m[38;2;31;10;0m█[0m[38;2;183;145;83m█[0m[38;2;174;134;75m█[0m[38;2;182;141;85m█[0m[38;2;184;143;87m█[0m[38;2;232;215;189m█[0m[38;2;226;214;190m█[0m[38;2;225;213;189m█[0m[38;2;224;214;189m██[0m[38;2;220;208;184m█[0m[38;2;224;212;188m█[0m[38;2;226;214;190m█[0m[38;2;35;25;13m█[0m[38;2;34;24;12m█[0m[38;2;50;49;44m█[0m[38;2;52;49;44m█[0m[38;2;53;50;43m█[0m[38;2;49;45;42m█[0m[38;2;64;63;58m█[0m[38;2;62;61;56m█[0m[38;2;54;51;46m█[0m");
$display("[38;2;41;41;39m█[0m[38;2;38;38;36m█[0m[38;2;39;39;37m█[0m[38;2;41;42;37m█[0m[38;2;83;100;110m█[0m[38;2;43;44;39m█[0m[38;2;42;41;39m█[0m[38;2;39;39;39m█[0m[38;2;46;45;40m█[0m[38;2;49;46;41m█[0m[38;2;47;44;39m█[0m[38;2;56;53;48m█[0m[38;2;56;51;45m█[0m[38;2;39;25;12m█[0m[38;2;33;20;11m█[0m[38;2;237;228;211m█[0m[38;2;226;212;186m█[0m[38;2;224;213;191m█[0m[38;2;223;213;186m█[0m[38;2;226;214;190m█[0m[38;2;223;211;187m██[0m[38;2;227;215;191m█[0m[38;2;224;212;188m█[0m[38;2;222;210;186m█[0m[38;2;226;215;193m█[0m[38;2;230;220;195m█[0m[38;2;221;211;186m█[0m[38;2;35;32;17m█[0m[38;2;154;105;100m█[0m[38;2;174;116;105m█[0m[38;2;164;104;94m█[0m[38;2;47;39;26m█[0m[38;2;167;110;99m█[0m[38;2;166;112;100m█[0m[38;2;173;113;103m█[0m[38;2;45;32;23m█[0m[38;2;255;248;231m█[0m[38;2;32;22;12m█[0m[38;2;245;237;218m█[0m[38;2;222;211;189m█[0m[38;2;222;210;186m█[0m[38;2;224;212;188m█[0m[38;2;232;220;196m█[0m[38;2;229;217;193m█[0m[38;2;225;213;189m██[0m[38;2;228;216;192m█[0m[38;2;233;221;197m█[0m[38;2;222;210;186m█[0m[38;2;226;214;190m█[0m[38;2;224;212;190m█[0m[38;2;223;213;188m█[0m[38;2;225;213;189m█[0m[38;2;224;212;188m█[0m[38;2;222;210;186m█[0m[38;2;229;218;196m█[0m[38;2;116;110;94m█[0m[38;2;36;23;14m█[0m[38;2;42;26;11m█[0m[38;2;41;27;14m█[0m[38;2;179;140;75m█[0m[38;2;178;137;83m█[0m[38;2;183;143;84m█[0m[38;2;188;148;89m█[0m[38;2;181;141;82m█[0m[38;2;180;139;83m█[0m[38;2;180;138;80m█[0m[38;2;183;141;83m█[0m[38;2;181;139;81m█[0m[38;2;184;144;85m█[0m[38;2;181;140;84m█[0m[38;2;187;147;88m█[0m[38;2;183;143;84m█[0m[38;2;187;147;88m█[0m[38;2;219;177;135m█[0m[38;2;36;27;10m█[0m[38;2;99;138;167m█[0m[38;2;34;21;12m█[0m[38;2;182;142;81m█[0m[38;2;179;138;82m█[0m[38;2;179;137;79m█[0m[38;2;181;139;81m█[0m[38;2;220;214;192m█[0m[38;2;224;212;188m█[0m[38;2;223;211;187m█[0m[38;2;224;212;188m█[0m[38;2;223;211;187m█[0m[38;2;224;212;188m█[0m[38;2;226;214;190m█[0m[38;2;224;212;188m█[0m[38;2;213;206;187m█[0m[38;2;33;21;9m█[0m[38;2;41;40;35m█[0m[38;2;38;38;36m█[0m[38;2;39;39;37m█[0m[38;2;35;35;33m█[0m[38;2;41;41;39m█[0m[38;2;48;47;43m█[0m[38;2;49;48;44m█[0m");
$display("[38;2;53;52;48m█[0m[38;2;50;49;45m█[0m[38;2;60;59;54m█[0m[38;2;48;45;40m█[0m[38;2;53;50;45m█[0m[38;2;66;75;80m█[0m[38;2;45;44;39m█[0m[38;2;48;47;42m█[0m[38;2;44;43;38m█[0m[38;2;52;49;44m█[0m[38;2;50;47;42m█[0m[38;2;53;50;43m█[0m[38;2;42;26;11m█[0m[38;2;38;26;14m█[0m[38;2;36;24;12m█[0m[38;2;38;26;14m█[0m[38;2;31;21;9m█[0m[38;2;224;215;200m█[0m[38;2;230;218;196m█[0m[38;2;226;216;191m█[0m[38;2;224;212;188m█[0m[38;2;229;217;193m█[0m[38;2;221;209;185m█[0m[38;2;224;214;189m█[0m[38;2;229;219;194m█[0m[38;2;229;217;193m█[0m[38;2;224;212;188m█[0m[38;2;226;214;190m█[0m[38;2;226;224;212m█[0m[38;2;47;33;24m█[0m[38;2;114;65;51m█[0m[38;2;169;109;101m█[0m[38;2;167;107;97m█[0m[38;2;174;116;105m█[0m[38;2;162;111;92m█[0m[38;2;45;32;23m█[0m[38;2;38;28;18m█[0m[38;2;227;215;191m█[0m[38;2;222;210;186m█[0m[38;2;226;214;190m█[0m[38;2;224;212;188m██[0m[38;2;228;216;192m█[0m[38;2;226;214;190m██[0m[38;2;224;212;188m█[0m[38;2;226;214;190m█[0m[38;2;223;211;187m█[0m[38;2;226;214;190m█[0m[38;2;228;216;192m█[0m[38;2;221;210;188m█[0m[38;2;7;0;0m█[0m[38;2;33;23;13m█[0m[38;2;36;24;8m█[0m[38;2;40;23;15m█[0m[38;2;33;20;11m█[0m[38;2;35;24;20m█[0m[38;2;177;141;81m█[0m[38;2;184;141;88m█[0m[38;2;194;147;95m█[0m[38;2;181;141;80m█[0m[38;2;179;139;80m███[0m[38;2;180;140;81m█[0m[38;2;186;146;87m█[0m[38;2;190;150;91m█[0m[38;2;189;147;89m██[0m[38;2;183;142;86m█[0m[38;2;179;137;79m█[0m[38;2;184;142;84m█[0m[38;2;183;141;83m██[0m[38;2;181;139;81m█[0m[38;2;154;118;56m█[0m[38;2;171;138;93m█[0m[38;2;5;1;2m█[0m[38;2;168;115;61m█[0m[38;2;149;113;55m█[0m[38;2;148;108;57m█[0m[38;2;151;109;61m█[0m[38;2;129;105;69m█[0m[38;2;35;25;16m█[0m[38;2;177;162;139m█[0m[38;2;184;169;146m█[0m[38;2;163;151;127m█[0m[38;2;177;165;141m█[0m[38;2;173;161;137m█[0m[38;2;161;146;123m█[0m[38;2;176;160;137m█[0m[38;2;20;6;0m█[0m[38;2;36;24;12m█[0m[38;2;41;42;37m█[0m[38;2;47;47;45m█[0m[38;2;49;48;44m█[0m[38;2;47;46;42m█[0m[38;2;53;52;47m██[0m[38;2;51;48;41m█[0m");
$display("[38;2;56;55;50m██[0m[38;2;53;50;41m█[0m[38;2;53;50;43m█[0m[38;2;47;44;39m█[0m[38;2;58;57;52m█[0m[38;2;49;50;44m█[0m[38;2;49;48;43m█[0m[38;2;49;49;41m█[0m[38;2;51;50;45m█[0m[38;2;38;24;13m█[0m[38;2;40;26;15m█[0m[38;2;255;255;243m█[0m[38;2;225;213;189m█[0m[38;2;228;216;192m██[0m[38;2;251;243;224m█[0m[38;2;39;25;12m█[0m[38;2;39;27;15m█[0m[38;2;38;25;16m█[0m[38;2;9;3;0m█[0m[38;2;234;219;196m█[0m[38;2;228;216;190m█[0m[38;2;222;215;189m█[0m[38;2;223;211;187m█[0m[38;2;224;213;191m██[0m[38;2;224;212;190m█[0m[38;2;228;216;192m█[0m[38;2;223;211;187m█[0m[38;2;228;218;193m█[0m[38;2;255;251;233m█[0m[38;2;23;15;4m█[0m[38;2;65;57;44m█[0m[38;2;255;245;223m█[0m[38;2;222;211;189m█[0m[38;2;220;210;185m█[0m[38;2;222;210;186m█[0m[38;2;224;212;188m█[0m[38;2;225;213;189m█[0m[38;2;229;217;193m█[0m[38;2;227;215;191m█[0m[38;2;226;214;190m█[0m[38;2;222;210;186m█[0m[38;2;224;212;186m█[0m[38;2;227;216;188m█[0m[38;2;228;216;190m█[0m[38;2;128;116;104m█[0m[38;2;35;23;11m█[0m[38;2;37;25;13m█[0m[38;2;32;19;10m█[0m[38;2;6;0;0m█[0m[38;2;223;211;187m█[0m[38;2;229;219;194m█[0m[38;2;223;211;187m█[0m[38;2;226;214;190m█[0m[38;2;171;142;100m█[0m[38;2;189;150;91m█[0m[38;2;180;137;86m█[0m[38;2;178;138;79m█[0m[38;2;181;141;82m█[0m[38;2;178;138;79m█[0m[38;2;181;141;80m█[0m[38;2;182;143;84m█[0m[38;2;184;143;87m█[0m[38;2;185;142;87m█[0m[38;2;186;146;87m█[0m[38;2;184;141;86m█[0m[38;2;175;136;81m█[0m[38;2;226;204;167m█[0m[38;2;229;214;191m█[0m[38;2;229;219;194m█[0m[38;2;181;166;145m█[0m[38;2;175;160;139m█[0m[38;2;170;155;134m█[0m[38;2;149;114;74m█[0m[38;2;168;130;83m█[0m[38;2;156;112;63m█[0m[38;2;153;113;64m█[0m[38;2;156;114;66m█[0m[38;2;144;112;63m█[0m[38;2;53;31;7m█[0m[38;2;34;25;10m█[0m[38;2;36;24;12m█[0m[38;2;97;84;68m█[0m[38;2;159;142;122m█[0m[38;2;175;157;135m█[0m[38;2;180;164;139m█[0m[38;2;176;159;139m█[0m[38;2;10;0;0m█[0m[38;2;38;25;16m█[0m[38;2;35;27;16m█[0m[38;2;40;44;45m█[0m[38;2;58;63;67m█[0m[38;2;65;74;79m█[0m[38;2;62;71;76m█[0m[38;2;65;74;79m█[0m[38;2;50;54;57m█[0m[38;2;55;52;47m█[0m[38;2;62;59;54m█[0m");
$display("[38;2;52;51;46m█[0m[38;2;51;50;45m█[0m[38;2;50;50;48m█[0m[38;2;81;82;84m█[0m[38;2;68;69;71m█[0m[38;2;69;70;72m█[0m[38;2;47;49;46m█[0m[38;2;46;45;40m█[0m[38;2;49;48;44m█[0m[38;2;38;25;16m█[0m[38;2;28;18;8m█[0m[38;2;226;216;191m█[0m[38;2;227;215;193m█[0m[38;2;215;207;184m█[0m[38;2;226;214;190m█[0m[38;2;227;215;191m█[0m[38;2;228;216;192m█[0m[38;2;226;214;190m█[0m[38;2;224;212;188m█[0m[38;2;231;223;202m█[0m[38;2;29;15;2m█[0m[38;2;34;24;14m█[0m[38;2;35;23;11m█[0m[38;2;32;20;8m█[0m[38;2;41;29;17m█[0m[38;2;11;0;0m█[0m[38;2;155;139;124m█[0m[38;2;169;151;129m█[0m[38;2;173;156;136m█[0m[38;2;183;166;146m█[0m[38;2;181;166;145m█[0m[38;2;184;169;148m█[0m[38;2;174;159;138m█[0m[38;2;176;161;140m██[0m[38;2;196;184;162m█[0m[38;2;176;161;140m█[0m[38;2;180;165;144m█[0m[38;2;178;163;142m██[0m[38;2;174;159;138m█[0m[38;2;180;165;144m█[0m[38;2;189;174;153m█[0m[38;2;178;163;142m█[0m[38;2;182;170;148m█[0m[38;2;210;199;181m█[0m[38;2;39;27;15m█[0m[38;2;33;20;11m█[0m[38;2;212;204;185m█[0m[38;2;223;213;186m█[0m[38;2;224;212;188m█[0m[38;2;226;214;190m█[0m[38;2;228;216;192m█[0m[38;2;223;211;187m██[0m[38;2;224;212;188m█[0m[38;2;223;211;187m█[0m[38;2;225;213;189m█[0m[38;2;233;216;198m█[0m[38;2;182;139;86m█[0m[38;2;177;141;81m█[0m[38;2;187;146;90m█[0m[38;2;177;137;78m█[0m[38;2;183;143;84m█[0m[38;2;186;149;97m█[0m[38;2;175;144;87m█[0m[38;2;150;142;123m█[0m[38;2;174;159;136m█[0m[38;2;180;165;142m█[0m[38;2;174;159;138m█[0m[38;2;178;163;142m█[0m[38;2;173;158;137m█[0m[38;2;179;164;143m█[0m[38;2;180;165;144m█[0m[38;2;174;159;138m█[0m[38;2;177;161;138m██[0m[38;2;175;160;141m█[0m[38;2;12;0;0m█[0m[38;2;45;32;24m█[0m[38;2;33;23;14m█[0m[38;2;35;23;11m█[0m[38;2;36;32;29m█[0m[38;2;28;23;17m█[0m[38;2;32;22;12m█[0m[38;2;31;21;11m█[0m[38;2;36;24;12m██[0m[38;2;34;24;14m█[0m[38;2;27;26;22m█[0m[38;2;32;36;39m█[0m[38;2;37;41;44m█[0m[38;2;32;36;37m█[0m[38;2;26;31;35m█[0m[38;2;67;76;81m█[0m[38;2;63;68;74m█[0m[38;2;60;69;76m█[0m[38;2;54;56;55m█[0m[38;2;54;51;46m█[0m[38;2;52;49;44m█[0m");
$display("[38;2;64;63;58m█[0m[38;2;66;65;60m█[0m[38;2;64;63;58m█[0m[38;2;53;52;47m█[0m[38;2;46;45;40m█[0m[38;2;50;49;44m█[0m[38;2;53;53;45m█[0m[38;2;46;47;41m█[0m[38;2;36;38;35m█[0m[38;2;34;21;12m█[0m[38;2;30;20;10m█[0m[38;2;225;211;185m█[0m[38;2;36;25;19m█[0m[38;2;211;202;185m█[0m[38;2;228;216;192m█[0m[38;2;227;215;191m█[0m[38;2;255;248;232m█[0m[38;2;226;215;193m█[0m[38;2;225;213;189m█[0m[38;2;222;210;186m█[0m[38;2;174;159;138m█[0m[38;2;187;172;151m█[0m[38;2;175;160;137m█[0m[38;2;178;162;139m█[0m[38;2;183;172;152m█[0m[38;2;38;25;16m█[0m[38;2;35;22;13m█[0m[38;2;36;24;12m█[0m[38;2;35;23;11m█[0m[38;2;36;24;12m█[0m[38;2;32;20;8m█[0m[38;2;32;22;12m█[0m[38;2;30;20;11m█[0m[38;2;37;25;13m█[0m[38;2;21;9;0m█[0m[38;2;69;57;43m█[0m[38;2;214;201;184m█[0m[38;2;184;171;152m█[0m[38;2;174;162;140m██[0m[38;2;166;154;132m█[0m[38;2;174;159;138m█[0m[38;2;176;163;144m█[0m[38;2;170;157;138m█[0m[38;2;41;27;16m█[0m[38;2;37;25;9m█[0m[38;2;208;197;175m█[0m[38;2;229;217;193m█[0m[38;2;225;215;188m█[0m[38;2;225;213;187m█[0m[38;2;230;218;194m█[0m[38;2;226;214;190m█[0m[38;2;227;215;191m█[0m[38;2;228;216;192m█[0m[38;2;225;213;189m██[0m[38;2;224;212;188m█[0m[38;2;222;210;186m█[0m[38;2;223;211;187m█[0m[38;2;228;211;183m█[0m[38;2;196;151;94m█[0m[38;2;187;146;90m█[0m[38;2;184;145;80m█[0m[38;2;179;143;81m█[0m[38;2;29;18;12m█[0m[38;2;38;26;14m█[0m[38;2;177;161;138m█[0m[38;2;173;159;133m█[0m[38;2;187;173;147m█[0m[38;2;190;175;152m█[0m[38;2;185;170;151m█[0m[38;2;58;46;32m█[0m[38;2;36;26;14m█[0m[38;2;36;26;16m█[0m[38;2;33;23;11m█[0m[38;2;33;23;13m█[0m[38;2;33;24;9m█[0m[38;2;33;21;9m█[0m[38;2;26;21;15m█[0m[38;2;28;35;41m█[0m[38;2;26;31;34m█[0m[38;2;31;35;38m█[0m[38;2;30;34;37m█[0m[38;2;35;39;42m█[0m[38;2;31;35;38m█[0m[38;2;36;40;43m█[0m[38;2;32;37;40m█[0m[38;2;33;37;38m█[0m[38;2;34;38;39m█[0m[38;2;31;35;36m█[0m[38;2;33;37;40m█[0m[38;2;62;71;76m█[0m[38;2;53;62;67m█[0m[38;2;58;67;72m█[0m[38;2;59;58;53m█[0m[38;2;55;52;47m█[0m[38;2;54;51;46m██[0m[38;2;57;56;51m█[0m[38;2;53;52;47m█[0m");
$display("[38;2;56;53;48m█[0m[38;2;53;50;45m██[0m[38;2;55;52;47m█[0m[38;2;49;46;41m█[0m[38;2;54;50;47m█[0m[38;2;34;35;37m█[0m[38;2;34;38;39m█[0m[38;2;29;33;34m█[0m[38;2;30;35;39m█[0m[38;2;37;25;13m█[0m[38;2;37;24;15m█[0m[38;2;35;25;15m█[0m[38;2;34;26;15m█[0m[38;2;150;146;134m█[0m[38;2;212;203;186m█[0m[38;2;37;25;13m█[0m[38;2;22;14;1m█[0m[38;2;11;1;0m█[0m[38;2;42;29;21m█[0m[38;2;33;23;11m█[0m[38;2;34;24;12m█[0m[38;2;33;23;11m█[0m[38;2;39;23;8m█[0m[38;2;37;23;12m█[0m[38;2;33;30;25m█[0m[38;2;34;39;42m█[0m[38;2;33;37;38m█[0m[38;2;34;38;39m█[0m[38;2;32;37;40m█[0m[38;2;31;35;36m█[0m[38;2;22;29;35m█[0m[38;2;38;42;43m█[0m[38;2;34;34;32m█[0m[38;2;33;26;18m█[0m[38;2;36;27;20m█[0m[38;2;36;24;12m█[0m[38;2;41;29;15m█[0m[38;2;38;24;11m█[0m[38;2;37;23;14m█[0m[38;2;40;26;17m█[0m[38;2;37;25;11m█[0m[38;2;36;22;13m█[0m[38;2;35;21;12m█[0m[38;2;34;22;10m█[0m[38;2;7;0;0m█[0m[38;2;226;214;192m█[0m[38;2;254;246;227m█[0m[38;2;33;24;15m█[0m[38;2;228;218;193m█[0m[38;2;229;217;193m█[0m[38;2;219;207;183m█[0m[38;2;255;249;232m█[0m[38;2;222;211;191m█[0m[38;2;224;212;186m█[0m[38;2;224;212;188m██[0m[38;2;227;215;191m█[0m[38;2;221;209;185m█[0m[38;2;224;214;187m█[0m[38;2;224;216;193m█[0m[38;2;23;0;0m█[0m[38;2;31;23;12m█[0m[38;2;35;23;7m█[0m[38;2;37;25;13m█[0m[38;2;37;24;15m█[0m[38;2;35;22;13m█[0m[38;2;37;25;13m█[0m[38;2;40;28;16m█[0m[38;2;35;21;10m█[0m[38;2;36;22;9m█[0m[38;2;32;22;12m█[0m[38;2;44;44;44m█[0m[38;2;29;33;34m█[0m[38;2;31;35;38m█[0m[38;2;25;30;33m█[0m[38;2;31;35;36m█[0m[38;2;30;35;38m█[0m[38;2;31;35;38m█[0m[38;2;32;36;39m█[0m[38;2;38;43;46m█[0m[38;2;34;40;40m█[0m[38;2;58;65;73m█[0m[38;2;57;66;71m█[0m[38;2;61;70;75m█[0m[38;2;56;65;70m█[0m[38;2;61;70;75m█[0m[38;2;62;71;76m█[0m[38;2;71;80;85m█[0m[38;2;63;72;77m█[0m[38;2;58;67;72m█[0m[38;2;57;66;73m█[0m[38;2;67;76;83m█[0m[38;2;65;74;81m█[0m[38;2;69;78;83m█[0m[38;2;66;74;77m█[0m[38;2;45;44;40m█[0m[38;2;53;50;45m█[0m[38;2;48;45;40m█[0m[38;2;51;48;43m█[0m");
$display("[38;2;48;47;42m█[0m[38;2;52;51;46m█[0m[38;2;53;52;47m█[0m[38;2;63;69;69m█[0m[38;2;61;68;74m█[0m[38;2;58;67;72m█[0m[38;2;63;70;76m█[0m[38;2;57;65;68m█[0m[38;2;34;39;43m█[0m[38;2;41;49;51m█[0m[38;2;36;40;41m█[0m[38;2;32;36;37m█[0m[38;2;36;41;45m█[0m[38;2;39;39;39m█[0m[38;2;39;36;31m█[0m[38;2;33;30;25m██[0m[38;2;33;32;27m█[0m[38;2;38;37;33m█[0m[38;2;30;32;31m█[0m[38;2;30;35;38m█[0m[38;2;31;36;40m█[0m[38;2;33;37;38m█[0m[38;2;31;35;38m█[0m[38;2;28;32;35m█[0m[38;2;33;37;40m██[0m[38;2;28;33;36m█[0m[38;2;33;37;40m█[0m[38;2;30;34;37m█[0m[38;2;33;37;40m█[0m[38;2;31;36;39m██[0m[38;2;35;39;42m█[0m[38;2;28;32;35m█[0m[38;2;35;39;42m█[0m[38;2;32;37;40m█[0m[38;2;29;34;37m██[0m[38;2;33;38;41m█[0m[38;2;29;34;37m█[0m[38;2;29;33;36m█[0m[38;2;33;37;40m█[0m[38;2;32;36;39m█[0m[38;2;34;22;10m█[0m[38;2;31;19;7m█[0m[38;2;127;117;105m█[0m[38;2;33;22;16m█[0m[38;2;73;65;46m█[0m[38;2;223;213;188m█[0m[38;2;226;214;190m█[0m[38;2;217;205;181m█[0m[38;2;35;21;8m█[0m[38;2;225;213;187m█[0m[38;2;222;212;187m█[0m[38;2;220;208;184m█[0m[38;2;215;208;182m█[0m[38;2;255;254;236m█[0m[38;2;31;19;7m█[0m[38;2;34;21;12m█[0m[38;2;34;24;12m█[0m[38;2;33;24;15m█[0m[38;2;25;35;37m█[0m[38;2;30;34;35m█[0m[38;2;32;36;37m█[0m[38;2;31;35;36m██[0m[38;2;29;33;36m█[0m[38;2;27;31;34m█[0m[38;2;33;37;40m█[0m[38;2;32;37;40m█[0m[38;2;28;33;36m█[0m[38;2;31;36;39m█[0m[38;2;30;35;38m█[0m[38;2;31;36;39m█[0m[38;2;55;62;68m█[0m[38;2;61;68;74m█[0m[38;2;55;62;68m█[0m[38;2;53;62;67m█[0m[38;2;51;60;65m█[0m[38;2;60;69;74m█[0m[38;2;59;68;73m█[0m[38;2;56;65;70m█[0m[38;2;62;71;76m█[0m[38;2;68;77;82m█[0m[38;2;58;67;72m█[0m[38;2;63;72;79m█[0m[38;2;67;75;78m█[0m[38;2;55;59;60m█[0m[38;2;51;52;47m█[0m[38;2;52;53;48m█[0m[38;2;49;46;39m█[0m[38;2;65;62;57m█[0m[38;2;53;50;45m█[0m[38;2;57;58;53m█[0m[38;2;48;47;42m█[0m[38;2;51;50;45m█[0m[38;2;48;47;42m█[0m[38;2;55;52;47m█[0m[38;2;54;51;46m█[0m");
$display("[38;2;47;46;41m█[0m[38;2;52;51;46m█[0m[38;2;49;48;43m█[0m[38;2;47;47;39m█[0m[38;2;54;62;64m█[0m[38;2;60;68;71m█[0m[38;2;58;65;71m█[0m[38;2;57;64;70m█[0m[38;2;62;69;75m█[0m[38;2;58;66;69m█[0m[38;2;57;65;68m█[0m[38;2;54;62;65m█[0m[38;2;36;41;44m█[0m[38;2;41;45;48m█[0m[38;2;35;39;42m█[0m[38;2;36;40;43m█[0m[38;2;31;35;38m██[0m[38;2;37;41;44m█[0m[38;2;34;38;41m█[0m[38;2;38;43;46m█[0m[38;2;37;41;42m█[0m[38;2;31;35;36m█[0m[38;2;37;41;44m█[0m[38;2;38;43;46m█[0m[38;2;34;38;41m█[0m[38;2;33;37;40m█[0m[38;2;34;39;42m█[0m[38;2;32;37;40m█[0m[38;2;27;32;35m█[0m[38;2;32;36;39m█[0m[38;2;31;35;38m█[0m[38;2;32;36;39m█[0m[38;2;36;41;44m█[0m[38;2;34;38;41m█[0m[38;2;37;41;44m█[0m[38;2;31;35;38m█[0m[38;2;28;33;36m█[0m[38;2;37;42;45m█[0m[38;2;27;32;35m██[0m[38;2;27;31;34m█[0m[38;2;32;36;39m█[0m[38;2;27;31;34m█[0m[38;2;28;34;32m█[0m[38;2;18;29;35m█[0m[38;2;34;25;18m█[0m[38;2;39;27;15m█[0m[38;2;33;23;14m█[0m[38;2;35;20;13m█[0m[38;2;34;24;14m█[0m[38;2;33;23;13m█[0m[38;2;39;26;17m█[0m[38;2;34;24;12m█[0m[38;2;31;21;11m█[0m[38;2;36;26;16m█[0m[38;2;33;26;10m█[0m[38;2;38;21;13m█[0m[38;2;37;36;34m█[0m[38;2;34;33;31m█[0m[38;2;35;40;44m█[0m[38;2;42;46;49m█[0m[38;2;30;35;38m█[0m[38;2;33;38;41m█[0m[38;2;31;36;39m█[0m[38;2;32;37;40m█[0m[38;2;28;33;36m█[0m[38;2;31;36;39m██[0m[38;2;35;39;42m█[0m[38;2;31;36;39m██[0m[38;2;29;34;37m█[0m[38;2;35;40;44m█[0m[38;2;32;36;37m█[0m[38;2;35;40;43m█[0m[38;2;73;82;87m█[0m[38;2;59;68;73m█[0m[38;2;60;69;74m█[0m[38;2;86;95;100m█[0m[38;2;93;98;102m██[0m[38;2;95;100;104m█[0m[38;2;87;95;98m█[0m[38;2;56;65;70m█[0m[38;2;63;72;77m█[0m[38;2;63;74;80m█[0m[38;2;66;76;78m█[0m[38;2;52;51;46m█[0m[38;2;54;51;46m█[0m[38;2;51;48;43m█[0m[38;2;43;44;39m█[0m[38;2;35;39;38m█[0m[38;2;33;37;36m█[0m[38;2;38;39;41m█[0m[38;2;39;41;40m█[0m[38;2;36;37;39m█[0m[38;2;39;41;40m█[0m[38;2;37;37;35m█[0m[38;2;34;34;32m█[0m");
$display("[38;2;50;49;44m█[0m[38;2;45;44;39m█[0m[38;2;48;47;42m█[0m[38;2;47;46;41m█[0m[38;2;45;44;39m█[0m[38;2;49;48;43m██[0m[38;2;48;47;42m█[0m[38;2;45;44;39m█[0m[38;2;54;53;48m█[0m[38;2;51;50;45m█[0m[38;2;48;47;42m█[0m[38;2;52;51;46m█[0m[38;2;57;61;62m█[0m[38;2;56;63;69m█[0m[38;2;55;62;68m█[0m[38;2;53;62;67m█[0m[38;2;56;65;70m█[0m[38;2;54;63;68m█[0m[38;2;64;73;78m█[0m[38;2;56;65;70m█[0m[38;2;58;67;72m█[0m[38;2;56;63;69m█[0m[38;2;51;60;65m█[0m[38;2;62;71;76m█[0m[38;2;54;63;68m█[0m[38;2;53;62;67m█[0m[38;2;58;67;72m█[0m[38;2;57;66;71m█[0m[38;2;36;41;45m█[0m[38;2;31;36;39m█[0m[38;2;34;39;42m█[0m[38;2;33;38;41m█[0m[38;2;39;43;46m█[0m[38;2;43;47;50m█[0m[38;2;38;42;45m█[0m[38;2;61;65;64m█[0m[38;2;49;53;54m██[0m[38;2;48;52;53m█[0m[38;2;49;54;57m█[0m[38;2;44;48;51m█[0m[38;2;37;42;45m█[0m[38;2;30;35;38m█[0m[38;2;34;39;42m█[0m[38;2;28;33;36m█[0m[38;2;34;39;42m█[0m[38;2;31;34;39m█[0m[38;2;31;35;38m█[0m[38;2;32;36;39m█[0m[38;2;35;39;42m██[0m[38;2;31;35;38m█[0m[38;2;28;32;35m█[0m[38;2;31;35;38m█[0m[38;2;31;36;39m██[0m[38;2;35;40;43m█[0m[38;2;33;37;40m█[0m[38;2;29;34;38m█[0m[38;2;35;40;44m█[0m[38;2;54;63;68m█[0m[38;2;55;62;68m█[0m[38;2;56;63;69m█[0m[38;2;60;67;73m█[0m[38;2;58;65;71m█[0m[38;2;54;63;68m█[0m[38;2;57;66;71m█[0m[38;2;58;67;72m█[0m[38;2;55;64;69m█[0m[38;2;56;65;72m█[0m[38;2;57;66;73m█[0m[38;2;55;64;71m██[0m[38;2;61;70;77m█[0m[38;2;67;76;83m█[0m[38;2;60;69;76m█[0m[38;2;76;85;90m█[0m[38;2;53;63;72m█[0m[38;2;72;85;91m█[0m[38;2;66;77;83m█[0m[38;2;63;74;80m█[0m[38;2;60;71;77m█[0m[38;2;64;75;79m█[0m[38;2;60;69;76m█[0m[38;2;65;74;79m█[0m[38;2;65;76;82m█[0m[38;2;65;72;78m█[0m[38;2;55;52;45m█[0m[38;2;51;50;45m█[0m[38;2;48;47;42m█[0m[38;2;55;52;47m█[0m[38;2;58;55;50m█[0m[38;2;53;50;45m█[0m[38;2;45;44;39m█[0m[38;2;41;41;39m█[0m[38;2;40;40;38m█[0m[38;2;33;35;32m█[0m[38;2;35;36;31m█[0m[38;2;43;44;39m█[0m");
$display("[38;2;36;36;36m█[0m[38;2;33;33;33m█[0m[38;2;34;36;35m█[0m[38;2;36;38;37m█[0m[38;2;34;36;35m█[0m[38;2;44;44;44m█[0m[38;2;34;34;34m█[0m[38;2;39;39;39m█[0m[38;2;38;38;36m█[0m[38;2;55;54;49m█[0m[38;2;51;50;45m█[0m[38;2;46;45;40m█[0m[38;2;53;52;47m█[0m[38;2;58;66;69m█[0m[38;2;58;67;72m█[0m[38;2;59;70;76m█[0m[38;2;59;67;70m█[0m[38;2;56;64;67m█[0m[38;2;60;68;71m█[0m[38;2;66;74;77m█[0m[38;2;68;76;79m█[0m[38;2;56;64;67m█[0m[38;2;60;68;71m█[0m[38;2;64;72;75m█[0m[38;2;58;66;69m█[0m[38;2;60;69;74m█[0m[38;2;61;70;75m█[0m[38;2;55;64;69m█[0m[38;2;67;72;76m█[0m[38;2;31;36;39m█[0m[38;2;33;37;40m█[0m[38;2;35;39;42m█[0m[38;2;34;38;41m█[0m[38;2;28;32;35m█[0m[38;2;29;33;36m█[0m[38;2;30;34;37m█[0m[38;2;32;36;37m██[0m[38;2;31;35;36m█[0m[38;2;52;57;60m█[0m[38;2;60;69;76m█[0m[38;2;65;74;79m█[0m[38;2;60;69;74m█[0m[38;2;61;70;75m█[0m[38;2;65;74;79m█[0m[38;2;53;62;67m█[0m[38;2;59;68;73m█[0m[38;2;62;71;76m█[0m[38;2;64;73;80m█[0m[38;2;60;69;76m█[0m[38;2;58;67;74m█[0m[38;2;66;75;82m█[0m[38;2;70;79;84m█[0m[38;2;58;67;74m█[0m[38;2;57;66;73m█[0m[38;2;58;67;72m█[0m[38;2;54;63;70m█[0m[38;2;67;76;83m█[0m[38;2;59;68;75m█[0m[38;2;55;64;69m█[0m[38;2;60;69;74m█[0m[38;2;59;68;73m█[0m[38;2;98;106;109m█[0m[38;2;87;95;98m█[0m[38;2;90;98;101m█[0m[38;2;91;99;102m█[0m[38;2;94;102;105m█[0m[38;2;58;67;72m█[0m[38;2;66;75;80m█[0m[38;2;64;73;80m█[0m[38;2;62;71;76m█[0m[38;2;50;51;53m█[0m[38;2;54;53;49m█[0m[38;2;51;50;45m█[0m[38;2;55;52;47m█[0m[38;2;53;52;48m██[0m[38;2;64;61;56m█[0m[38;2;58;55;50m█[0m[38;2;55;52;47m█[0m[38;2;81;91;100m█[0m[38;2;54;51;46m█[0m[38;2;60;59;54m█[0m[38;2;56;53;48m█[0m[38;2;53;52;47m█[0m[38;2;55;54;49m█[0m[38;2;52;52;44m█[0m[38;2;51;48;43m█[0m[38;2;50;47;42m█[0m[38;2;57;54;49m█[0m[38;2;50;47;42m█[0m[38;2;71;70;66m█[0m[38;2;72;71;67m█[0m[38;2;71;70;66m█[0m[38;2;67;66;61m█[0m[38;2;49;46;41m█[0m[38;2;55;52;47m██[0m[38;2;57;54;49m█[0m[38;2;62;59;54m█[0m");
$display("[38;2;51;50;45m█[0m[38;2;50;49;45m█[0m[38;2;50;49;44m█[0m[38;2;44;45;40m█[0m[38;2;40;40;38m█[0m[38;2;33;33;33m█[0m[38;2;34;34;34m█[0m[38;2;36;36;36m█[0m[38;2;37;37;35m█[0m[38;2;41;40;36m█[0m[38;2;49;46;41m█[0m[38;2;48;47;42m█[0m[38;2;47;46;41m█[0m[38;2;49;48;43m█[0m[38;2;45;44;39m█[0m[38;2;51;50;45m█[0m[38;2;51;48;43m█[0m[38;2;53;50;45m█[0m[38;2;51;48;43m█[0m[38;2;50;49;44m█[0m[38;2;53;50;45m█[0m[38;2;52;49;44m█[0m[38;2;54;51;46m█[0m[38;2;53;50;41m█[0m[38;2;69;75;75m█[0m[38;2;57;66;71m█[0m[38;2;63;72;79m█[0m[38;2;59;68;73m█[0m[38;2;61;70;77m█[0m[38;2;58;67;74m█[0m[38;2;60;69;74m█[0m[38;2;58;67;72m█[0m[38;2;59;68;73m█[0m[38;2;64;73;80m█[0m[38;2;63;72;79m█[0m[38;2;57;66;73m█[0m[38;2;59;68;75m█[0m[38;2;60;69;74m█[0m[38;2;64;73;78m█[0m[38;2;58;65;71m█[0m[38;2;64;71;77m█[0m[38;2;71;78;84m█[0m[38;2;65;74;79m█[0m[38;2;63;70;76m█[0m[38;2;58;67;72m█[0m[38;2;61;70;75m█[0m[38;2;67;76;81m█[0m[38;2;61;69;72m█[0m[38;2;64;72;75m█[0m[38;2;66;74;77m█[0m[38;2;69;77;80m█[0m[38;2;66;74;77m█[0m[38;2;61;68;74m█[0m[38;2;63;72;77m█[0m[38;2;67;76;81m█[0m[38;2;61;70;75m█[0m[38;2;59;68;75m█[0m[38;2;56;65;72m█[0m[38;2;66;75;80m█[0m[38;2;62;71;78m█[0m[38;2;63;72;79m██[0m[38;2;57;66;71m█[0m[38;2;61;70;75m█[0m[38;2;60;69;74m█[0m[38;2;58;67;72m█[0m[38;2;66;74;77m█[0m[38;2;58;64;64m█[0m[38;2;49;49;47m█[0m[38;2;52;51;47m█[0m[38;2;52;49;44m██[0m[38;2;58;57;52m█[0m[38;2;47;44;39m█[0m[38;2;52;49;44m█[0m[38;2;53;50;45m█[0m[38;2;56;53;48m█[0m[38;2;50;47;42m█[0m[38;2;51;48;43m█[0m[38;2;53;50;45m█[0m[38;2;65;62;55m█[0m[38;2;93;107;116m█[0m[38;2;52;49;42m█[0m[38;2;47;46;41m█[0m[38;2;52;51;47m█[0m[38;2;50;49;45m█[0m[38;2;47;46;42m█[0m[38;2;50;49;44m█[0m[38;2;53;52;47m█[0m[38;2;54;51;46m█[0m[38;2;52;49;44m█[0m[38;2;46;45;40m█[0m[38;2;51;50;45m█[0m[38;2;43;42;37m█[0m[38;2;42;41;36m█[0m[38;2;51;50;45m█[0m[38;2;46;45;40m█[0m[38;2;55;54;49m█[0m[38;2;51;50;45m██[0m");
$display("[38;2;55;54;49m█[0m[38;2;49;48;43m█[0m[38;2;55;54;50m█[0m[38;2;39;39;37m█[0m[38;2;36;36;34m█[0m[38;2;33;35;34m█[0m[38;2;37;39;38m█[0m[38;2;38;40;39m█[0m[38;2;40;40;38m█[0m[38;2;40;40;40m█[0m[38;2;33;33;33m█[0m[38;2;36;38;37m█[0m[38;2;43;43;41m█[0m[38;2;48;47;42m█[0m[38;2;50;49;44m█[0m[38;2;55;54;49m█[0m[38;2;53;52;47m█[0m[38;2;51;50;45m█[0m[38;2;46;45;40m█[0m[38;2;50;49;44m██[0m[38;2;49;48;43m█[0m[38;2;50;49;44m█[0m[38;2;52;51;46m█[0m[38;2;53;50;45m█[0m[38;2;40;42;41m█[0m[38;2;59;67;69m█[0m[38;2;53;64;70m█[0m[38;2;58;69;75m█[0m[38;2;63;70;78m█[0m[38;2;63;72;77m█[0m[38;2;59;68;75m█[0m[38;2;63;72;79m█[0m[38;2;67;76;83m█[0m[38;2;74;84;93m█[0m[38;2;64;73;78m█[0m[38;2;69;78;85m█[0m[38;2;63;72;77m█[0m[38;2;64;73;78m█[0m[38;2;56;65;70m█[0m[38;2;64;73;78m█[0m[38;2;70;79;84m█[0m[38;2;71;80;85m█[0m[38;2;56;65;70m█[0m[38;2;56;65;72m█[0m[38;2;58;71;79m█[0m[38;2;58;67;72m█[0m[38;2;62;67;70m█[0m[38;2;51;48;43m█[0m[38;2;53;50;45m██[0m[38;2;50;47;42m██[0m[38;2;58;55;50m█[0m[38;2;52;49;44m█[0m[38;2;58;55;50m█[0m[38;2;51;48;43m█[0m[38;2;53;50;45m█[0m[38;2;60;57;52m█[0m[38;2;55;52;47m█[0m[38;2;47;44;39m█[0m[38;2;62;59;54m█[0m[38;2;48;47;42m█[0m[38;2;49;48;43m█[0m[38;2;54;51;46m█[0m[38;2;52;49;44m█[0m[38;2;63;60;55m█[0m[38;2;53;50;45m█[0m[38;2;51;48;43m██[0m[38;2;54;53;48m█[0m[38;2;48;47;42m█[0m[38;2;51;50;46m█[0m[38;2;39;41;40m█[0m[38;2;37;39;38m█[0m[38;2;38;40;39m██[0m[38;2;36;38;37m█[0m[38;2;36;38;35m█[0m[38;2;58;57;55m█[0m[38;2;44;43;38m█[0m[38;2;52;49;44m█[0m[38;2;74;82;85m█[0m[38;2;49;46;41m█[0m[38;2;48;45;40m█[0m[38;2;54;51;46m█[0m[38;2;46;45;40m█[0m[38;2;49;46;41m█[0m[38;2;51;48;43m█[0m[38;2;56;53;48m█[0m[38;2;59;56;51m█[0m[38;2;55;54;50m█[0m[38;2;40;39;35m█[0m[38;2;39;38;34m█[0m[38;2;43;42;38m█[0m[38;2;46;45;41m█[0m[38;2;44;43;39m█[0m[38;2;49;48;44m█[0m[38;2;48;47;42m██[0m");
$display("[38;2;52;51;46m█[0m[38;2;47;46;41m█[0m[38;2;49;48;43m█[0m[38;2;55;52;47m█[0m[38;2;52;49;44m█[0m[38;2;49;48;43m█[0m[38;2;47;44;39m█[0m[38;2;50;47;42m█[0m[38;2;63;60;55m█[0m[38;2;51;50;45m█[0m[38;2;61;60;55m█[0m[38;2;55;52;47m█[0m[38;2;53;50;45m█[0m[38;2;54;53;48m█[0m[38;2;49;48;43m█[0m[38;2;54;53;48m█[0m[38;2;40;40;38m█[0m[38;2;38;38;36m██[0m[38;2;39;39;37m█[0m[38;2;36;36;34m█[0m[38;2;42;42;40m█[0m[38;2;57;56;52m█[0m[38;2;50;49;44m█[0m[38;2;52;51;46m██[0m[38;2;49;48;43m█[0m[38;2;52;51;46m█[0m[38;2;51;50;45m█[0m[38;2;55;54;49m█[0m[38;2;56;56;48m█[0m[38;2;57;58;52m█[0m[38;2;53;52;48m█[0m[38;2;45;44;39m█[0m[38;2;55;56;50m█[0m[38;2;52;57;53m█[0m[38;2;41;45;44m█[0m[38;2;53;52;48m█[0m[38;2;50;49;45m█[0m[38;2;49;50;44m█[0m[38;2;47;48;42m█[0m[38;2;50;49;45m█[0m[38;2;48;48;40m█[0m[38;2;56;52;49m█[0m[38;2;53;50;45m█[0m[38;2;50;47;42m█[0m[38;2;51;48;43m█[0m[38;2;52;49;44m██[0m[38;2;56;53;48m█[0m[38;2;50;49;44m█[0m[38;2;51;50;45m█[0m[38;2;55;52;47m█[0m[38;2;50;49;44m█[0m[38;2;47;46;41m█[0m[38;2;57;56;52m█[0m[38;2;37;37;35m█[0m[38;2;37;39;38m█[0m[38;2;36;38;37m██[0m[38;2;38;40;39m█[0m[38;2;35;37;36m█[0m[38;2;42;41;36m█[0m[38;2;48;47;42m█[0m[38;2;52;51;46m█[0m[38;2;51;50;45m█[0m[38;2;43;44;39m█[0m[38;2;41;43;42m█[0m[38;2;34;36;35m█[0m[38;2;34;34;34m█[0m[38;2;32;32;32m█[0m[38;2;33;33;33m█[0m[38;2;31;33;32m█[0m[38;2;36;38;37m█[0m[38;2;33;35;34m█[0m[38;2;34;36;35m█[0m[38;2;38;40;39m█[0m[38;2;35;37;36m█[0m[38;2;43;45;44m█[0m[38;2;37;39;38m█[0m[38;2;35;35;35m█[0m[38;2;35;37;36m█[0m[38;2;32;34;33m█[0m[38;2;35;37;36m█[0m[38;2;33;35;34m█[0m[38;2;39;41;40m█[0m[38;2;37;37;37m█[0m[38;2;45;44;39m█[0m[38;2;50;49;44m█[0m[38;2;52;49;44m█[0m[38;2;49;46;41m█[0m[38;2;49;48;43m█[0m[38;2;52;51;46m█[0m[38;2;50;49;44m██[0m[38;2;54;53;48m█[0m[38;2;47;46;41m█[0m[38;2;49;48;43m█[0m[38;2;50;49;44m█[0m[38;2;51;50;45m█[0m");
$display("[38;2;50;49;44m█[0m[38;2;48;47;42m█[0m[38;2;45;44;39m█[0m[38;2;50;49;44m█[0m[38;2;53;52;47m█[0m[38;2;54;53;48m█[0m[38;2;48;47;42m█[0m[38;2;53;52;47m█[0m[38;2;51;50;45m█[0m[38;2;50;51;43m█[0m[38;2;38;38;36m█[0m[38;2;33;35;34m█[0m[38;2;36;38;37m█[0m[38;2;35;37;36m█[0m[38;2;29;30;32m█[0m[38;2;31;35;34m█[0m[38;2;35;37;36m█[0m[38;2;44;44;44m█[0m[38;2;36;36;36m█[0m[38;2;36;38;37m█[0m[38;2;37;39;38m█[0m[38;2;31;33;32m█[0m[38;2;45;47;42m█[0m[38;2;47;46;41m█[0m[38;2;50;49;44m█[0m[38;2;48;47;42m█[0m[38;2;53;52;47m█[0m[38;2;51;50;45m█[0m[38;2;46;45;40m█[0m[38;2;48;47;42m█[0m[38;2;45;44;39m█[0m[38;2;47;44;39m█[0m[38;2;50;47;42m█[0m[38;2;51;50;45m█[0m[38;2;47;46;41m█[0m[38;2;48;47;42m█[0m[38;2;46;43;38m█[0m[38;2;108;105;100m█[0m[38;2;53;50;45m█[0m[38;2;53;52;47m█[0m[38;2;54;53;48m█[0m[38;2;49;46;41m█[0m[38;2;51;48;43m█[0m[38;2;54;51;46m█[0m[38;2;50;49;44m█[0m[38;2;49;48;43m█[0m[38;2;50;49;44m██[0m[38;2;49;48;43m█[0m[38;2;54;53;48m█[0m[38;2;49;48;43m█[0m[38;2;36;40;41m█[0m[38;2;37;39;36m█[0m[38;2;36;38;37m█[0m[38;2;34;36;35m██[0m[38;2;35;37;36m█[0m[38;2;37;39;38m█[0m[38;2;33;35;34m██[0m[38;2;41;43;42m█[0m[38;2;40;42;39m█[0m[38;2;50;46;43m█[0m[38;2;48;47;42m█[0m[38;2;49;46;41m█[0m[38;2;53;50;45m█[0m[38;2;55;52;47m█[0m[38;2;57;54;49m█[0m[38;2;49;46;41m█[0m[38;2;47;46;41m█[0m[38;2;52;49;44m█[0m[38;2;56;53;48m█[0m[38;2;50;49;44m█[0m[38;2;41;43;40m█[0m[38;2;33;35;32m█[0m[38;2;34;36;35m█[0m[38;2;36;38;37m█[0m[38;2;38;40;39m█[0m[38;2;33;35;34m█[0m[38;2;32;34;33m█[0m[38;2;38;40;39m█[0m[38;2;37;39;38m█[0m[38;2;36;38;37m█[0m[38;2;32;34;33m█[0m[38;2;36;38;37m█[0m[38;2;32;34;33m█[0m[38;2;35;37;36m█[0m[38;2;36;36;34m█[0m[38;2;34;34;32m█[0m[38;2;37;37;37m██[0m[38;2;39;41;38m█[0m[38;2;42;41;36m█[0m[38;2;49;48;43m█[0m[38;2;52;51;46m█[0m[38;2;51;48;43m█[0m[38;2;56;53;48m█[0m[38;2;50;47;42m█[0m[38;2;51;48;43m█[0m[38;2;58;55;50m█[0m");
$display("[38;2;41;42;37m█[0m[38;2;43;44;39m█[0m[38;2;39;40;35m█[0m[38;2;41;41;39m██[0m[38;2;43;42;38m█[0m[38;2;45;44;40m█[0m[38;2;52;51;47m█[0m[38;2;45;44;39m█[0m[38;2;50;49;44m█[0m[38;2;47;46;41m█[0m[38;2;50;49;44m█[0m[38;2;51;50;45m█[0m[38;2;37;37;35m█[0m[38;2;31;31;29m█[0m[38;2;37;37;35m█[0m[38;2;34;34;32m█[0m[38;2;34;36;35m█[0m[38;2;37;39;38m█[0m[38;2;35;39;38m█[0m[38;2;35;37;36m█[0m[38;2;37;39;38m█[0m[38;2;39;39;37m█[0m[38;2;45;44;39m█[0m[38;2;52;51;46m██[0m[38;2;54;53;48m█[0m[38;2;50;49;44m█[0m[38;2;42;43;38m█[0m[38;2;40;40;38m█[0m[38;2;32;32;30m█[0m[38;2;39;39;39m█[0m[38;2;36;36;36m█[0m[38;2;50;49;44m█[0m[38;2;49;48;43m██[0m[38;2;53;52;47m█[0m[38;2;54;46;35m█[0m[38;2;69;78;83m█[0m[38;2;50;49;44m█[0m[38;2;47;46;41m█[0m[38;2;51;48;43m█[0m[38;2;52;51;46m█[0m[38;2;50;49;44m█[0m[38;2;51;50;45m█[0m[38;2;53;50;45m█[0m[38;2;56;53;48m█[0m[38;2;52;51;46m█[0m[38;2;50;47;42m█[0m[38;2;55;52;47m█[0m[38;2;51;48;43m█[0m[38;2;44;41;36m█[0m[38;2;52;51;46m█[0m[38;2;57;54;49m█[0m[38;2;50;47;42m█[0m[38;2;47;46;41m█[0m[38;2;51;48;43m█[0m[38;2;52;49;44m█[0m[38;2;50;47;42m█[0m[38;2;50;49;44m█[0m[38;2;40;41;36m█[0m[38;2;44;44;42m█[0m[38;2;47;44;39m█[0m[38;2;48;47;42m██[0m[38;2;49;48;43m███[0m[38;2;46;45;40m█[0m[38;2;54;53;48m█[0m[38;2;52;51;46m█[0m[38;2;48;47;42m█[0m[38;2;49;48;43m█[0m[38;2;53;52;47m█[0m[38;2;49;48;43m█[0m[38;2;55;52;47m█[0m[38;2;54;51;46m█[0m[38;2;51;50;45m█[0m[38;2;50;49;45m██[0m[38;2;52;49;44m█[0m[38;2;46;45;40m█[0m[38;2;48;47;42m█[0m[38;2;59;58;53m█[0m[38;2;52;49;44m██[0m[38;2;50;47;42m█[0m[38;2;45;44;39m█[0m[38;2;47;46;41m█[0m[38;2;46;45;40m█[0m[38;2;47;46;41m█[0m[38;2;52;51;46m█[0m[38;2;50;49;44m█[0m[38;2;47;46;42m█[0m[38;2;46;45;40m█[0m[38;2;44;43;39m██[0m[38;2;42;43;38m█[0m[38;2;43;42;38m█[0m[38;2;42;41;37m█[0m");
$display("[38;2;43;44;39m█[0m[38;2;44;45;40m█[0m[38;2;42;42;40m█[0m[38;2;44;44;42m██[0m[38;2;46;46;44m█[0m[38;2;44;45;40m█[0m[38;2;43;44;39m█[0m[38;2;46;45;41m█[0m[38;2;44;43;39m█[0m[38;2;48;47;43m█[0m[38;2;46;45;40m█[0m[38;2;50;49;44m█[0m[38;2;49;48;43m█[0m[38;2;46;45;40m█[0m[38;2;50;49;44m█[0m[38;2;53;50;45m█[0m[38;2;54;53;48m█[0m[38;2;60;59;54m█[0m[38;2;54;53;48m█[0m[38;2;50;49;44m█[0m[38;2;56;55;50m█[0m[38;2;51;50;45m█[0m[38;2;46;45;40m█[0m[38;2;54;53;48m█[0m[38;2;48;47;42m█[0m[38;2;52;51;46m█[0m[38;2;48;47;42m█[0m[38;2;51;48;43m█[0m[38;2;48;45;40m█[0m[38;2;44;43;38m█[0m[38;2;52;51;46m█[0m[38;2;51;50;45m█[0m[38;2;48;47;42m█[0m[38;2;50;49;44m█[0m[38;2;52;51;46m██[0m[38;2;53;50;45m█[0m[38;2;49;46;41m█[0m[38;2;48;47;42m█[0m[38;2;49;48;43m█[0m[38;2;48;47;42m█[0m[38;2;50;49;44m█[0m[38;2;49;48;43m█[0m[38;2;51;50;45m███[0m[38;2;45;44;39m█[0m[38;2;50;49;44m█[0m[38;2;54;53;48m█[0m[38;2;49;46;41m█[0m[38;2;50;47;42m█[0m[38;2;48;47;42m█[0m[38;2;51;48;43m█[0m[38;2;54;51;46m█[0m[38;2;48;47;42m█[0m[38;2;56;55;50m█[0m[38;2;54;53;48m█[0m[38;2;52;49;44m█[0m[38;2;52;51;46m█[0m[38;2;55;54;49m█[0m[38;2;51;50;45m█[0m[38;2;49;48;43m█[0m[38;2;52;51;46m█[0m[38;2;46;45;40m█[0m[38;2;50;49;44m█[0m[38;2;55;54;49m█[0m[38;2;50;49;44m█[0m[38;2;46;45;40m█[0m[38;2;43;42;38m█[0m[38;2;44;45;40m█[0m[38;2;43;44;39m█[0m[38;2;50;49;44m█[0m[38;2;51;50;45m█[0m[38;2;54;53;48m█[0m[38;2;46;45;40m█[0m[38;2;44;43;38m█[0m[38;2;49;48;43m██[0m[38;2;51;50;45m█[0m[38;2;57;56;51m█[0m[38;2;55;54;49m█[0m[38;2;54;53;48m█[0m[38;2;47;46;41m█[0m[38;2;50;49;44m█[0m[38;2;48;47;42m█[0m[38;2;46;45;41m█[0m[38;2;47;46;42m█[0m[38;2;46;45;41m█[0m[38;2;48;47;43m█[0m[38;2;50;49;45m█[0m[38;2;51;50;46m█[0m[38;2;46;45;41m█[0m[38;2;41;40;36m█[0m[38;2;41;41;39m█[0m[38;2;42;41;37m█[0m[38;2;43;42;38m█[0m[38;2;44;45;40m█[0m[38;2;40;39;35m█[0m[38;2;47;46;42m█[0m");    
    $display("\n");
    $display("                         \033[31m\033[5m █████ █████ █████ █████ █████ \033[0m");
    $display("                         \033[31m\033[5m █     █   █ █   █ █   █ █   █ \033[0m");
    $display("                         \033[31m\033[5m █████ █████ █████ █   █ █████ \033[0m");
    $display("                         \033[31m\033[5m █     █  █  █  █  █   █ █  █  \033[0m");
    $display("                         \033[31m\033[5m █████ █   █ █   █ █████ █   █ \033[0m");
    $display("\n");
end endtask      



task display_pass; begin
    $display("[38;2;209;198;123m█[0m[38;2;189;193;139m█[0m[38;2;184;191;135m█[0m[38;2;191;195;136m█[0m[38;2;197;194;132m█[0m[38;2;197;195;130m█[0m[38;2;195;192;133m█[0m[38;2;195;196;134m█[0m[38;2;196;197;136m█[0m[38;2;193;197;135m█[0m[38;2;179;194;143m█[0m[38;2;179;193;143m█[0m[38;2;171;189;145m█[0m[38;2;154;189;151m█[0m[38;2;156;188;150m█[0m[38;2;175;194;148m█[0m[38;2;163;189;148m█[0m[38;2;157;188;154m█[0m[38;2;143;187;159m█[0m[38;2;142;188;164m█[0m[38;2;129;180;164m█[0m[38;2;120;176;167m█[0m[38;2;120;178;169m█[0m[38;2;119;182;170m█[0m[38;2;120;180;169m█[0m[38;2;137;182;158m█[0m[38;2;143;183;156m█[0m[38;2;137;180;156m█[0m[38;2;124;175;161m█[0m[38;2;130;182;167m█[0m[38;2;127;181;167m█[0m[38;2;125;179;168m█[0m[38;2;120;179;170m█[0m[38;2;114;181;173m█[0m[38;2;105;176;174m█[0m[38;2;98;170;173m█[0m[38;2;86;167;173m█[0m[38;2;83;169;180m█[0m[38;2;80;167;180m█[0m[38;2;63;159;179m█[0m[38;2;62;160;182m█[0m[38;2;63;161;183m█[0m[38;2;61;158;180m█[0m[38;2;58;156;180m█[0m[38;2;60;154;179m█[0m[38;2;56;153;183m█[0m[38;2;56;154;181m█[0m[38;2;58;152;181m█[0m[38;2;54;153;180m█[0m[38;2;58;153;182m█[0m[38;2;60;158;184m█[0m[38;2;53;152;179m█[0m[38;2;58;157;180m█[0m[38;2;54;152;181m█[0m[38;2;57;155;182m█[0m[38;2;53;154;179m█[0m[38;2;54;152;183m█[0m[38;2;54;153;183m█[0m[38;2;47;149;178m█[0m[38;2;45;151;186m█[0m[38;2;39;142;181m█[0m[38;2;40;148;184m█[0m[38;2;32;143;179m█[0m[38;2;30;136;180m█[0m[38;2;31;143;183m█[0m[38;2;30;140;182m█[0m[38;2;27;137;180m█[0m[38;2;29;140;184m█[0m[38;2;30;139;182m█[0m[38;2;27;137;182m█[0m[38;2;28;140;182m█[0m[38;2;30;139;184m█[0m[38;2;29;143;186m█[0m[38;2;30;140;184m█[0m[38;2;26;136;182m█[0m[38;2;26;136;181m█[0m[38;2;25;137;185m█[0m[38;2;27;139;183m█[0m[38;2;27;140;185m█[0m[38;2;29;137;184m█[0m[38;2;30;140;184m█[0m[38;2;26;136;181m█[0m[38;2;24;136;182m█[0m[38;2;26;138;184m█[0m[38;2;24;139;182m█[0m[38;2;25;136;185m█[0m[38;2;22;135;180m█[0m[38;2;24;137;181m█[0m[38;2;26;137;185m█[0m[38;2;23;136;182m█[0m[38;2;24;140;184m█[0m[38;2;25;139;183m█[0m[38;2;27;139;186m█[0m[38;2;26;139;186m█[0m[38;2;26;138;184m█[0m[38;2;26;142;187m█[0m[38;2;24;137;184m█[0m[38;2;18;134;179m█[0m[38;2;27;141;187m█[0m[38;2;28;141;186m█[0m");
$display("[38;2;217;203;121m█[0m[38;2;219;202;121m█[0m[38;2;199;197;130m█[0m[38;2;202;197;129m█[0m[38;2;205;198;125m█[0m[38;2;210;198;122m█[0m[38;2;219;199;123m█[0m[38;2;215;199;123m█[0m[38;2;212;199;127m█[0m[38;2;215;203;127m█[0m[38;2;205;197;131m█[0m[38;2;200;199;134m█[0m[38;2;194;195;138m█[0m[38;2;187;193;136m█[0m[38;2;192;196;134m█[0m[38;2;195;197;134m█[0m[38;2;182;194;139m█[0m[38;2;174;193;148m█[0m[38;2;162;190;151m█[0m[38;2;163;191;160m█[0m[38;2;151;184;153m█[0m[38;2;154;184;150m█[0m[38;2;155;188;155m█[0m[38;2;170;190;147m█[0m[38;2;171;193;147m█[0m[38;2;158;189;154m█[0m[38;2;152;184;156m█[0m[38;2;157;192;161m█[0m[38;2;155;190;160m█[0m[38;2;147;186;156m█[0m[38;2;138;178;156m█[0m[38;2;132;185;165m█[0m[38;2;124;182;167m█[0m[38;2;99;173;175m█[0m[38;2;100;172;173m█[0m[38;2;97;171;171m█[0m[38;2;89;168;176m█[0m[38;2;86;171;177m█[0m[38;2;85;166;174m█[0m[38;2;81;165;174m█[0m[38;2;87;171;181m█[0m[38;2;77;163;176m█[0m[38;2;76;164;182m█[0m[38;2;73;163;178m█[0m[38;2;69;161;180m█[0m[38;2;71;162;178m█[0m[38;2;69;159;176m█[0m[38;2;66;159;181m█[0m[38;2;65;158;180m█[0m[38;2;64;160;181m█[0m[38;2;66;158;176m█[0m[38;2;66;158;180m█[0m[38;2;63;158;183m█[0m[38;2;59;159;183m█[0m[38;2;57;155;181m█[0m[38;2;51;154;183m█[0m[38;2;45;150;181m█[0m[38;2;41;151;184m█[0m[38;2;38;144;180m█[0m[38;2;37;147;187m█[0m[38;2;32;143;182m█[0m[38;2;31;144;185m█[0m[38;2;32;142;186m█[0m[38;2;29;141;187m█[0m[38;2;29;142;184m█[0m[38;2;29;143;184m█[0m[38;2;29;141;184m█[0m[38;2;32;144;187m█[0m[38;2;29;143;186m█[0m[38;2;30;144;189m█[0m[38;2;26;142;182m█[0m[38;2;29;146;189m█[0m[38;2;27;142;183m█[0m[38;2;32;144;185m█[0m[38;2;30;144;187m█[0m[38;2;25;140;183m█[0m[38;2;31;143;185m█[0m[38;2;32;146;185m█[0m[38;2;30;146;187m█[0m[38;2;26;142;182m█[0m[38;2;35;150;189m█[0m[38;2;27;142;185m█[0m[38;2;29;144;187m█[0m[38;2;28;143;186m█[0m[38;2;27;147;185m█[0m[38;2;28;143;187m█[0m[38;2;25;140;184m█[0m[38;2;26;143;185m█[0m[38;2;29;147;187m█[0m[38;2;27;144;188m█[0m[38;2;34;152;190m█[0m[38;2;31;147;189m█[0m[38;2;26;143;184m█[0m[38;2;29;144;188m█[0m[38;2;26;141;186m█[0m[38;2;28;145;188m█[0m[38;2;29;147;192m█[0m[38;2;27;145;185m█[0m[38;2;25;143;184m█[0m[38;2;27;144;189m█[0m");
$display("[38;2;226;203;119m█[0m[38;2;229;202;117m█[0m[38;2;224;200;114m█[0m[38;2;221;202;121m█[0m[38;2;217;198;118m█[0m[38;2;228;204;116m█[0m[38;2;229;204;113m█[0m[38;2;233;205;112m█[0m[38;2;237;207;115m█[0m[38;2;239;209;119m█[0m[38;2;226;202;117m█[0m[38;2;221;199;118m█[0m[38;2;224;204;121m█[0m[38;2;220;203;120m█[0m[38;2;223;204;120m█[0m[38;2;219;204;123m█[0m[38;2;204;196;126m█[0m[38;2;192;197;136m█[0m[38;2;186;195;141m█[0m[38;2;189;196;140m█[0m[38;2;187;193;135m█[0m[38;2;200;199;136m█[0m[38;2;192;199;138m█[0m[38;2;191;196;141m█[0m[38;2;181;195;143m█[0m[38;2;179;196;144m█[0m[38;2;180;194;146m█[0m[38;2;172;195;152m█[0m[38;2;163;190;148m█[0m[38;2;143;187;161m█[0m[38;2;134;185;163m█[0m[38;2;131;183;165m█[0m[38;2;114;178;167m█[0m[38;2;112;176;168m█[0m[38;2;114;178;169m█[0m[38;2;122;181;169m█[0m[38;2;118;179;169m█[0m[38;2;102;169;165m█[0m[38;2;107;173;168m█[0m[38;2;114;179;167m█[0m[38;2;106;172;168m█[0m[38;2;99;175;173m█[0m[38;2;89;166;168m█[0m[38;2;90;169;175m█[0m[38;2;87;169;178m█[0m[38;2;87;170;176m█[0m[38;2;78;163;175m█[0m[38;2;82;170;181m█[0m[38;2;77;167;179m█[0m[38;2;71;160;179m█[0m[38;2;61;160;178m█[0m[38;2;57;157;186m█[0m[38;2;51;157;186m█[0m[38;2;45;154;185m█[0m[38;2;38;151;181m█[0m[38;2;36;148;184m█[0m[38;2;39;149;186m█[0m[38;2;35;151;184m█[0m[38;2;38;153;187m█[0m[38;2;34;147;184m█[0m[38;2;35;147;186m█[0m[38;2;37;150;186m█[0m[38;2;37;149;187m█[0m[38;2;35;150;186m█[0m[38;2;35;144;185m█[0m[38;2;33;147;184m█[0m[38;2;31;149;184m█[0m[38;2;39;151;190m█[0m[38;2;37;149;184m█[0m[38;2;32;146;186m█[0m[38;2;33;149;185m█[0m[38;2;35;151;186m█[0m[38;2;43;155;191m█[0m[38;2;33;148;182m█[0m[38;2;38;152;187m█[0m[38;2;37;152;185m█[0m[38;2;38;152;190m█[0m[38;2;38;154;190m█[0m[38;2;35;149;187m█[0m[38;2;29;144;184m█[0m[38;2;34;150;188m█[0m[38;2;29;146;184m█[0m[38;2;31;149;186m█[0m[38;2;35;151;190m█[0m[38;2;27;146;184m█[0m[38;2;28;144;186m█[0m[38;2;27;144;189m█[0m[38;2;26;143;182m█[0m[38;2;32;149;189m█[0m[38;2;27;144;185m█[0m[38;2;26;144;187m█[0m[38;2;28;147;189m█[0m[38;2;26;145;189m█[0m[38;2;25;145;188m█[0m[38;2;31;149;192m█[0m[38;2;32;151;190m█[0m[38;2;28;147;189m█[0m[38;2;27;145;188m█[0m[38;2;26;146;186m█[0m[38;2;32;152;191m█[0m");
$display("[38;2;225;204;119m█[0m[38;2;237;204;113m█[0m[38;2;239;208;111m█[0m[38;2;238;205;110m█[0m[38;2;231;201;109m█[0m[38;2;236;209;112m█[0m[38;2;243;207;107m█[0m[38;2;250;210;95m█[0m[38;2;250;207;92m█[0m[38;2;251;212;97m█[0m[38;2;252;210;94m█[0m[38;2;250;209;99m█[0m[38;2;246;206;104m█[0m[38;2;245;208;105m█[0m[38;2;238;209;111m█[0m[38;2;229;206;119m█[0m[38;2;221;203;118m█[0m[38;2;214;201;125m█[0m[38;2;217;204;126m█[0m[38;2;219;204;122m█[0m[38;2;215;199;125m█[0m[38;2;209;200;131m█[0m[38;2;199;198;131m█[0m[38;2;198;202;134m█[0m[38;2;190;197;139m█[0m[38;2;191;195;141m█[0m[38;2;168;191;152m█[0m[38;2;158;190;153m█[0m[38;2;154;185;151m█[0m[38;2;152;192;160m█[0m[38;2;145;189;157m█[0m[38;2;141;184;158m█[0m[38;2;146;187;161m█[0m[38;2;140;184;160m█[0m[38;2;141;186;160m█[0m[38;2;142;184;159m█[0m[38;2;130;181;162m█[0m[38;2;120;179;163m█[0m[38;2;120;177;166m█[0m[38;2;117;179;169m█[0m[38;2;111;177;170m█[0m[38;2;110;177;170m█[0m[38;2;104;174;176m█[0m[38;2;91;174;177m█[0m[38;2;83;170;183m█[0m[38;2;72;166;183m█[0m[38;2;73;168;184m█[0m[38;2;62;166;189m█[0m[38;2;53;160;188m█[0m[38;2;52;158;187m█[0m[38;2;48;158;187m█[0m[38;2;47;157;187m█[0m[38;2;50;159;189m█[0m[38;2;46;156;187m█[0m[38;2;53;166;197m█[0m[38;2;47;159;191m█[0m[38;2;47;155;189m█[0m[38;2;44;152;183m█[0m[38;2;45;154;190m█[0m[38;2;44;152;185m█[0m[38;2;46;157;187m█[0m[38;2;39;151;184m█[0m[38;2;44;155;187m█[0m[38;2;45;155;185m█[0m[38;2;44;152;183m█[0m[38;2;48;159;189m█[0m[38;2;51;159;187m█[0m[38;2;49;158;188m█[0m[38;2;49;160;188m█[0m[38;2;45;157;188m█[0m[38;2;46;157;189m█[0m[38;2;46;156;190m█[0m[38;2;43;157;190m█[0m[38;2;43;157;185m█[0m[38;2;41;154;187m█[0m[38;2;42;156;189m█[0m[38;2;41;157;195m█[0m[38;2;44;156;189m█[0m[38;2;34;152;189m█[0m[38;2;45;163;196m█[0m[38;2;35;152;186m█[0m[38;2;44;162;195m█[0m[38;2;30;149;187m█[0m[38;2;33;150;188m█[0m[38;2;35;155;187m█[0m[38;2;40;159;198m█[0m[38;2;31;151;188m█[0m[38;2;30;151;190m█[0m[38;2;32;149;188m█[0m[38;2;31;151;189m█[0m[38;2;27;147;186m█[0m[38;2;29;150;191m█[0m[38;2;30;151;191m█[0m[38;2;30;152;190m█[0m[38;2;26;149;191m█[0m[38;2;27;147;189m█[0m[38;2;32;154;194m█[0m[38;2;26;147;188m█[0m[38;2;27;149;190m█[0m[38;2;31;152;189m█[0m");
$display("[38;2;217;201;122m█[0m[38;2;227;202;118m█[0m[38;2;238;203;106m█[0m[38;2;251;210;102m█[0m[38;2;254;213;97m█[0m[38;2;253;212;94m█[0m[38;2;255;229;121m█[0m[38;2;254;227;120m█[0m[38;2;255;228;124m█[0m[38;2;254;227;117m█[0m[38;2;254;226;122m█[0m[38;2;255;228;123m█[0m[38;2;254;227;124m█[0m[38;2;253;216;96m█[0m[38;2;253;212;95m█[0m[38;2;249;209;98m█[0m[38;2;240;208;110m█[0m[38;2;244;211;115m█[0m[38;2;239;208;116m█[0m[38;2;227;204;120m█[0m[38;2;225;206;121m█[0m[38;2;213;205;125m█[0m[38;2;205;204;135m█[0m[38;2;181;197;139m█[0m[38;2;175;196;144m█[0m[38;2;175;196;149m█[0m[38;2;174;194;145m█[0m[38;2;170;193;150m█[0m[38;2;172;193;149m█[0m[38;2;174;194;149m█[0m[38;2;167;191;149m█[0m[38;2;162;190;149m█[0m[38;2;155;190;153m█[0m[38;2;149;189;156m█[0m[38;2;147;192;162m█[0m[38;2;136;186;160m█[0m[38;2;130;185;165m█[0m[38;2;113;181;171m█[0m[38;2;113;179;173m█[0m[38;2;107;175;178m█[0m[38;2;90;174;176m█[0m[38;2;78;169;180m█[0m[38;2;73;168;185m█[0m[38;2;64;168;181m█[0m[38;2;66;164;182m█[0m[38;2;66;165;183m█[0m[38;2;65;167;186m█[0m[38;2;66;166;189m█[0m[38;2;62;165;185m█[0m[38;2;56;164;187m█[0m[38;2;56;164;189m█[0m[38;2;58;161;187m█[0m[38;2;58;165;183m█[0m[38;2;57;160;186m█[0m[38;2;61;163;183m█[0m[38;2;61;160;188m█[0m[38;2;67;165;184m█[0m[38;2;63;163;183m█[0m[38;2;66;164;184m█[0m[38;2;68;166;186m█[0m[38;2;59;160;186m█[0m[38;2;56;160;188m█[0m[38;2;58;162;184m█[0m[38;2;51;160;187m█[0m[38;2;50;160;188m█[0m[38;2;53;164;193m█[0m[38;2;48;159;188m█[0m[38;2;45;157;192m█[0m[38;2;48;160;186m█[0m[38;2;45;157;190m█[0m[38;2;49;160;188m█[0m[38;2;43;155;188m█[0m[38;2;45;160;195m█[0m[38;2;37;156;190m█[0m[38;2;43;157;191m█[0m[38;2;51;165;199m█[0m[38;2;35;154;192m█[0m[38;2;36;158;195m█[0m[38;2;36;153;194m█[0m[38;2;28;151;189m█[0m[38;2;34;154;191m█[0m[38;2;30;153;193m█[0m[38;2;33;154;192m█[0m[38;2;32;152;192m█[0m[38;2;33;154;191m█[0m[38;2;31;154;193m█[0m[38;2;31;155;192m█[0m[38;2;38;157;193m█[0m[38;2;33;155;194m█[0m[38;2;32;154;190m█[0m[38;2;35;160;196m█[0m[38;2;34;159;195m█[0m[38;2;32;154;193m█[0m[38;2;31;155;193m█[0m[38;2;38;165;202m█[0m[38;2;32;154;193m█[0m[38;2;30;153;192m█[0m[38;2;28;153;192m█[0m[38;2;28;157;194m█[0m[38;2;36;163;201m█[0m");
$display("[38;2;228;206;116m█[0m[38;2;234;205;113m█[0m[38;2;249;209;96m█[0m[38;2;254;212;95m█[0m[38;2;253;227;127m█[0m[38;2;253;226;122m█[0m[38;2;255;229;127m█[0m[38;2;255;229;130m█[0m[38;2;252;230;134m█[0m[38;2;253;231;134m█[0m[38;2;254;230;137m█[0m[38;2;254;230;133m█[0m[38;2;255;231;134m█[0m[38;2;253;229;127m█[0m[38;2;254;231;127m█[0m[38;2;251;220;104m█[0m[38;2;254;217;99m█[0m[38;2;247;210;100m█[0m[38;2;240;208;113m█[0m[38;2;229;206;119m█[0m[38;2;216;204;123m█[0m[38;2;208;201;128m█[0m[38;2;204;203;135m█[0m[38;2;201;202;132m█[0m[38;2;207;203;134m█[0m[38;2;201;198;131m█[0m[38;2;200;200;135m█[0m[38;2;186;198;138m█[0m[38;2;181;196;142m█[0m[38;2;169;194;148m█[0m[38;2;162;192;151m█[0m[38;2;158;190;156m█[0m[38;2;150;190;153m█[0m[38;2;144;188;161m█[0m[38;2;134;188;165m█[0m[38;2;119;184;171m█[0m[38;2;109;183;175m█[0m[38;2;92;180;185m█[0m[38;2;89;177;182m█[0m[38;2;83;174;182m█[0m[38;2;79;170;181m█[0m[38;2;76;173;183m█[0m[38;2;85;175;187m█[0m[38;2;84;174;181m█[0m[38;2;88;173;181m█[0m[38;2;88;177;185m█[0m[38;2;88;175;183m█[0m[38;2;89;177;183m█[0m[38;2;84;173;183m█[0m[38;2;84;177;185m█[0m[38;2;78;171;183m█[0m[38;2;78;170;186m█[0m[38;2;78;170;181m█[0m[38;2;71;165;182m█[0m[38;2;68;168;186m█[0m[38;2;63;165;187m█[0m[38;2;64;164;184m█[0m[38;2;63;168;186m█[0m[38;2;63;164;191m█[0m[38;2;60;164;186m█[0m[38;2;54;161;189m█[0m[38;2;53;162;190m█[0m[38;2;49;162;188m█[0m[38;2;50;159;189m█[0m[38;2;49;163;190m█[0m[38;2;44;160;193m█[0m[38;2;44;161;192m█[0m[38;2;42;158;189m█[0m[38;2;36;157;188m█[0m[38;2;37;157;193m█[0m[38;2;37;159;194m█[0m[38;2;35;156;194m█[0m[38;2;33;155;191m█[0m[38;2;32;155;192m█[0m[38;2;34;156;192m█[0m[38;2;31;154;191m█[0m[38;2;37;159;198m█[0m[38;2;32;156;194m█[0m[38;2;33;159;196m█[0m[38;2;30;153;190m█[0m[38;2;31;158;195m█[0m[38;2;31;153;191m█[0m[38;2;35;158;195m█[0m[38;2;34;155;194m█[0m[38;2;39;162;195m█[0m[38;2;163;208;200m█[0m[38;2;195;217;201m█[0m[38;2;231;228;203m█[0m[38;2;236;228;200m█[0m[38;2;233;228;203m█[0m[38;2;224;225;198m█[0m[38;2;219;221;200m█[0m[38;2;139;200;209m█[0m[38;2;36;167;208m█[0m[38;2;37;162;199m█[0m[38;2;30;156;192m█[0m[38;2;30;155;194m█[0m[38;2;29;155;195m█[0m[38;2;27;155;192m█[0m[38;2;34;161;197m█[0m");
$display("[38;2;236;208;112m█[0m[38;2;249;211;100m█[0m[38;2;255;210;90m█[0m[38;2;255;228;124m█[0m[38;2;253;228;124m█[0m[38;2;252;228;129m█[0m[38;2;254;230;132m█[0m[38;2;253;233;145m█[0m[38;2;255;233;144m█[0m[38;2;254;233;145m█[0m[38;2;254;232;149m█[0m[38;2;254;233;142m█[0m[38;2;254;231;135m█[0m[38;2;255;233;135m█[0m[38;2;253;234;131m█[0m[38;2;255;230;129m█[0m[38;2;255;229;116m█[0m[38;2;254;214;98m█[0m[38;2;248;214;107m█[0m[38;2;240;209;109m█[0m[38;2;234;208;115m█[0m[38;2;226;206;114m█[0m[38;2;225;208;124m█[0m[38;2;215;206;127m█[0m[38;2;207;202;131m█[0m[38;2;194;197;133m█[0m[38;2;186;197;142m█[0m[38;2;176;195;145m█[0m[38;2;166;195;153m█[0m[38;2;152;192;160m█[0m[38;2;149;192;160m█[0m[38;2;137;186;159m█[0m[38;2;131;187;166m█[0m[38;2;131;185;167m█[0m[38;2;135;187;167m█[0m[38;2;133;189;168m█[0m[38;2;124;184;166m█[0m[38;2;120;184;168m█[0m[38;2;119;185;175m█[0m[38;2;109;180;174m█[0m[38;2;111;184;178m█[0m[38;2;107;181;175m█[0m[38;2;109;186;183m█[0m[38;2;98;182;183m█[0m[38;2;98;175;175m█[0m[38;2;101;183;181m█[0m[38;2;88;173;177m█[0m[38;2;88;177;182m█[0m[38;2;87;177;182m█[0m[38;2;83;172;180m█[0m[38;2;79;175;183m█[0m[38;2;72;170;187m█[0m[38;2;69;172;191m█[0m[38;2;61;167;191m█[0m[38;2;54;165;188m█[0m[38;2;52;165;191m█[0m[38;2;49;162;190m█[0m[38;2;40;162;192m█[0m[38;2;35;155;191m█[0m[38;2;41;158;192m█[0m[38;2;39;156;192m█[0m[38;2;35;158;192m█[0m[38;2;28;155;188m█[0m[38;2;32;154;191m█[0m[38;2;34;158;194m█[0m[38;2;32;156;192m█[0m[38;2;36;156;193m█[0m[38;2;37;161;196m█[0m[38;2;37;161;195m█[0m[38;2;33;154;190m█[0m[38;2;34;158;194m█[0m[38;2;33;156;195m█[0m[38;2;32;156;194m█[0m[38;2;31;158;192m█[0m[38;2;31;156;197m█[0m[38;2;32;158;197m█[0m[38;2;30;157;196m█[0m[38;2;32;158;195m█[0m[38;2;35;160;194m█[0m[38;2;28;155;192m█[0m[38;2;42;167;204m█[0m[38;2;34;162;200m█[0m[38;2;35;164;204m█[0m[38;2;208;222;202m█[0m[38;2;230;226;199m█[0m[38;2;237;230;199m█[0m[38;2;241;232;202m█[0m[38;2;241;232;199m█[0m[38;2;240;230;201m█[0m[38;2;239;232;202m█[0m[38;2;234;230;201m█[0m[38;2;226;226;201m█[0m[38;2;211;221;200m█[0m[38;2;212;222;201m█[0m[38;2;177;209;195m█[0m[38;2;36;164;199m█[0m[38;2;30;159;194m█[0m[38;2;34;161;197m█[0m[38;2;33;158;199m█[0m[38;2;30;154;190m█[0m");
$display("[38;2;240;209;112m█[0m[38;2;253;209;97m█[0m[38;2;254;226;122m█[0m[38;2;254;227;121m█[0m[38;2;254;229;129m█[0m[38;2;255;231;129m█[0m[38;2;253;233;139m█[0m[38;2;253;231;140m█[0m[38;2;252;233;149m█[0m[38;2;254;234;149m█[0m[38;2;254;232;143m██[0m[38;2;255;234;143m█[0m[38;2;255;234;137m█[0m[38;2;255;232;129m█[0m[38;2;255;231;125m█[0m[38;2;254;231;124m█[0m[38;2;255;218;96m█[0m[38;2;252;215;100m█[0m[38;2;241;212;110m█[0m[38;2;234;209;120m█[0m[38;2;217;202;125m█[0m[38;2;208;206;134m█[0m[38;2;192;203;139m█[0m[38;2;184;198;143m█[0m[38;2;175;199;152m█[0m[38;2;167;194;156m█[0m[38;2;164;195;156m█[0m[38;2;165;197;159m█[0m[38;2;151;192;163m█[0m[38;2;151;194;163m█[0m[38;2;152;195;164m█[0m[38;2;145;189;156m█[0m[38;2;154;198;162m█[0m[38;2;150;194;163m█[0m[38;2;140;190;164m█[0m[38;2;144;191;163m█[0m[38;2;131;188;167m█[0m[38;2;125;185;171m█[0m[38;2;118;183;171m█[0m[38;2;117;186;177m█[0m[38;2;106;182;180m█[0m[38;2;96;179;183m█[0m[38;2;83;178;185m█[0m[38;2;73;173;187m█[0m[38;2;67;172;191m█[0m[38;2;55;169;190m█[0m[38;2;50;166;194m█[0m[38;2;51;168;194m█[0m[38;2;43;164;194m█[0m[38;2;51;172;200m█[0m[38;2;40;164;197m█[0m[38;2;42;164;198m█[0m[38;2;39;167;196m█[0m[38;2;42;165;200m█[0m[38;2;39;161;193m█[0m[38;2;37;160;194m█[0m[38;2;36;161;197m█[0m[38;2;36;162;197m█[0m[38;2;34;158;193m█[0m[38;2;36;159;194m█[0m[38;2;39;162;194m█[0m[38;2;37;165;197m█[0m[38;2;34;162;201m█[0m[38;2;30;154;193m█[0m[38;2;30;157;197m█[0m[38;2;29;158;194m█[0m[38;2;34;161;198m█[0m[38;2;34;160;199m█[0m[38;2;32;158;195m█[0m[38;2;29;156;195m█[0m[38;2;31;158;195m█[0m[38;2;39;164;201m█[0m[38;2;31;161;196m█[0m[38;2;36;164;201m█[0m[38;2;33;159;198m█[0m[38;2;34;162;200m█[0m[38;2;32;160;196m█[0m[38;2;33;163;197m█[0m[38;2;33;162;198m█[0m[38;2;35;165;198m█[0m[38;2;38;171;213m█[0m[38;2;221;228;206m█[0m[38;2;241;233;202m█[0m[38;2;239;230;201m█[0m[38;2;240;231;201m█[0m[38;2;241;232;199m█[0m[38;2;235;231;199m█[0m[38;2;226;228;204m█[0m[38;2;223;225;198m█[0m[38;2;221;227;202m█[0m[38;2;179;216;204m█[0m[38;2;167;213;208m█[0m[38;2;178;218;205m█[0m[38;2;183;213;204m█[0m[38;2;152;206;208m█[0m[38;2;31;159;198m█[0m[38;2;34;162;193m█[0m[38;2;36;165;200m█[0m[38;2;35;164;201m█[0m");
$display("[38;2;235;206;108m█[0m[38;2;254;209;96m█[0m[38;2;252;228;122m█[0m[38;2;254;227;118m█[0m[38;2;255;229;123m█[0m[38;2;254;231;129m█[0m[38;2;253;231;138m█[0m[38;2;253;233;140m█[0m[38;2;253;235;148m█[0m[38;2;253;233;145m█[0m[38;2;255;234;144m█[0m[38;2;252;231;146m█[0m[38;2;255;232;144m█[0m[38;2;254;234;138m█[0m[38;2;254;232;128m█[0m[38;2;253;233;129m█[0m[38;2;253;229;121m█[0m[38;2;253;215;93m█[0m[38;2;248;212;104m█[0m[38;2;233;208;120m█[0m[38;2;222;208;128m█[0m[38;2;207;206;136m█[0m[38;2;195;201;138m█[0m[38;2;185;198;141m█[0m[38;2;180;202;152m█[0m[38;2;171;196;152m█[0m[38;2;168;194;154m█[0m[38;2;163;196;156m█[0m[38;2;156;194;161m█[0m[38;2;140;190;163m█[0m[38;2;135;191;168m█[0m[38;2;127;190;174m█[0m[38;2;118;184;177m█[0m[38;2;105;182;177m█[0m[38;2;104;182;177m█[0m[38;2;95;180;181m█[0m[38;2;90;181;185m█[0m[38;2;82;180;187m█[0m[38;2;76;177;187m█[0m[38;2;76;180;195m█[0m[38;2;66;173;189m█[0m[38;2;67;179;194m█[0m[38;2;62;172;193m█[0m[38;2;58;169;192m█[0m[38;2;57;174;194m█[0m[38;2;54;174;199m█[0m[38;2;55;174;199m█[0m[38;2;45;165;194m█[0m[38;2;45;166;199m█[0m[38;2;44;164;195m█[0m[38;2;46;169;199m█[0m[38;2;43;166;198m█[0m[38;2;35;162;193m█[0m[38;2;42;166;198m█[0m[38;2;40;167;197m█[0m[38;2;43;169;199m█[0m[38;2;43;167;199m█[0m[38;2;38;165;198m█[0m[38;2;37;164;197m█[0m[38;2;39;165;198m█[0m[38;2;34;164;198m█[0m[38;2;35;162;196m█[0m[38;2;35;165;199m█[0m[38;2;41;168;201m█[0m[38;2;35;164;197m█[0m[38;2;37;166;200m█[0m[38;2;36;166;198m█[0m[38;2;34;164;196m█[0m[38;2;34;164;198m█[0m[38;2;37;166;201m█[0m[38;2;33;162;196m█[0m[38;2;34;165;200m█[0m[38;2;38;167;203m█[0m[38;2;34;161;199m█[0m[38;2;31;162;198m█[0m[38;2;38;169;204m█[0m[38;2;40;170;206m█[0m[38;2;56;175;202m█[0m[38;2;67;182;207m█[0m[38;2;42;170;198m█[0m[38;2;43;174;204m█[0m[38;2;109;188;198m█[0m[38;2;224;227;201m█[0m[38;2;226;227;199m█[0m[38;2;229;227;198m█[0m[38;2;236;231;202m█[0m[38;2;221;226;203m█[0m[38;2;198;220;202m█[0m[38;2;188;217;204m█[0m[38;2;187;220;207m█[0m[38;2;169;213;205m█[0m[38;2;164;216;212m█[0m[38;2;160;213;208m█[0m[38;2;152;210;208m█[0m[38;2;157;211;209m█[0m[38;2;151;207;205m█[0m[38;2;35;166;200m█[0m[38;2;35;158;196m█[0m[38;2;78;177;198m█[0m[38;2;87;182;200m█[0m");
$display("[38;2;243;211;109m█[0m[38;2;250;209;99m█[0m[38;2;254;215;94m█[0m[38;2;255;231;125m█[0m[38;2;255;230;122m█[0m[38;2;254;231;130m█[0m[38;2;255;231;134m█[0m[38;2;253;230;136m█[0m[38;2;255;232;140m█[0m[38;2;253;231;138m█[0m[38;2;254;233;141m███[0m[38;2;255;228;126m█[0m[38;2;253;232;125m█[0m[38;2;254;232;126m█[0m[38;2;254;231;126m█[0m[38;2;252;216;97m█[0m[38;2;250;214;108m█[0m[38;2;237;208;114m█[0m[38;2;233;211;122m█[0m[38;2;222;206;126m█[0m[38;2;215;206;131m█[0m[38;2;196;203;136m█[0m[38;2;188;200;145m█[0m[38;2;180;199;148m█[0m[38;2;173;199;157m█[0m[38;2;160;196;157m█[0m[38;2;149;196;165m█[0m[38;2;133;193;174m█[0m[38;2;128;193;173m█[0m[38;2;121;188;176m█[0m[38;2;110;186;180m█[0m[38;2;104;186;188m█[0m[38;2;94;183;188m█[0m[38;2;94;183;187m█[0m[38;2;91;185;191m█[0m[38;2;78;180;193m█[0m[38;2;74;178;196m█[0m[38;2;70;178;192m█[0m[38;2;64;175;195m█[0m[38;2;63;175;196m█[0m[38;2;62;173;194m█[0m[38;2;59;175;195m█[0m[38;2;59;174;198m█[0m[38;2;53;172;195m█[0m[38;2;49;170;194m█[0m[38;2;53;171;198m█[0m[38;2;48;172;200m█[0m[38;2;48;169;198m█[0m[38;2;46;170;196m█[0m[38;2;50;169;201m█[0m[38;2;46;170;199m█[0m[38;2;43;170;198m█[0m[38;2;49;174;200m█[0m[38;2;44;171;199m█[0m[38;2;45;169;196m█[0m[38;2;48;173;203m█[0m[38;2;45;173;202m█[0m[38;2;47;172;203m█[0m[38;2;41;171;200m█[0m[38;2;44;169;199m█[0m[38;2;40;171;198m█[0m[38;2;39;168;200m█[0m[38;2;41;169;199m█[0m[38;2;36;163;198m█[0m[38;2;33;166;200m█[0m[38;2;38;168;202m█[0m[38;2;40;167;201m█[0m[38;2;33;166;198m█[0m[38;2;31;162;196m█[0m[38;2;37;169;202m█[0m[38;2;38;170;202m█[0m[38;2;37;169;199m█[0m[38;2;46;174;210m█[0m[38;2;205;224;206m█[0m[38;2;221;228;205m█[0m[38;2;233;229;203m█[0m[38;2;231;231;203m█[0m[38;2;221;228;202m█[0m[38;2;203;223;205m█[0m[38;2;205;221;202m█[0m[38;2;193;221;205m█[0m[38;2;204;223;202m█[0m[38;2;206;221;204m█[0m[38;2;209;224;206m█[0m[38;2;177;217;205m█[0m[38;2;167;217;211m█[0m[38;2;156;210;205m█[0m[38;2;145;210;205m█[0m[38;2;149;208;207m█[0m[38;2;138;203;205m█[0m[38;2;139;203;206m█[0m[38;2;143;206;206m█[0m[38;2;145;204;207m█[0m[38;2;143;205;206m█[0m[38;2;136;199;200m█[0m[38;2;140;201;203m█[0m[38;2;147;200;198m█[0m[38;2;139;198;200m█[0m");
$display("[38;2;218;202;117m█[0m[38;2;237;209;115m█[0m[38;2;253;209;90m█[0m[38;2;255;224;111m█[0m[38;2;254;227;118m█[0m[38;2;255;230;125m█[0m[38;2;255;226;117m█[0m[38;2;255;230;129m█[0m[38;2;254;228;124m█[0m[38;2;253;232;126m█[0m[38;2;255;229;124m█[0m[38;2;254;229;125m█[0m[38;2;251;232;134m█[0m[38;2;253;231;131m█[0m[38;2;254;232;128m█[0m[38;2;255;231;123m█[0m[38;2;254;219;99m█[0m[38;2;247;212;103m█[0m[38;2;231;210;116m█[0m[38;2;227;208;121m█[0m[38;2;226;209;127m█[0m[38;2;220;209;130m█[0m[38;2;212;206;133m██[0m[38;2;208;206;137m█[0m[38;2;194;202;140m█[0m[38;2;194;204;144m█[0m[38;2;184;205;154m█[0m[38;2;169;200;157m█[0m[38;2;157;200;168m█[0m[38;2;138;194;169m█[0m[38;2;136;192;169m█[0m[38;2;135;194;178m█[0m[38;2;125;190;177m█[0m[38;2;124;191;178m█[0m[38;2;118;188;179m█[0m[38;2;113;191;182m█[0m[38;2;108;189;182m█[0m[38;2;89;181;186m█[0m[38;2;80;181;186m█[0m[38;2;81;183;195m█[0m[38;2;66;176;194m█[0m[38;2;57;172;198m█[0m[38;2;59;176;199m█[0m[38;2;64;175;202m█[0m[38;2;49;170;198m█[0m[38;2;49;170;199m█[0m[38;2;52;176;202m█[0m[38;2;40;171;201m█[0m[38;2;43;169;199m█[0m[38;2;41;170;196m█[0m[38;2;43;172;202m█[0m[38;2;39;169;201m█[0m[38;2;41;170;198m█[0m[38;2;37;169;200m█[0m[38;2;41;171;201m█[0m[38;2;42;171;204m█[0m[38;2;40;168;203m█[0m[38;2;38;168;201m█[0m[38;2;36;166;201m█[0m[38;2;39;170;201m█[0m[38;2;33;167;200m█[0m[38;2;36;170;199m█[0m[38;2;43;170;203m█[0m[38;2;37;168;201m█[0m[38;2;38;169;202m█[0m[38;2;42;169;201m█[0m[38;2;51;178;211m█[0m[38;2;40;171;207m█[0m[38;2;43;173;204m█[0m[38;2;40;173;202m█[0m[38;2;43;174;205m█[0m[38;2;46;173;206m█[0m[38;2;50;177;204m█[0m[38;2;143;201;199m█[0m[38;2;222;229;210m█[0m[38;2;231;230;204m█[0m[38;2;227;229;204m█[0m[38;2;219;229;201m█[0m[38;2;204;228;208m█[0m[38;2;166;214;207m█[0m[38;2;171;216;206m█[0m[38;2;158;214;211m█[0m[38;2;165;211;202m█[0m[38;2;178;217;210m█[0m[38;2;160;212;203m█[0m[38;2;172;213;208m█[0m[38;2;138;207;208m█[0m[38;2;137;208;209m█[0m[38;2;135;206;208m█[0m[38;2;134;202;205m█[0m[38;2;133;203;209m█[0m[38;2;140;207;206m█[0m[38;2;133;201;205m█[0m[38;2;135;198;205m█[0m[38;2;135;199;204m█[0m[38;2;132;199;204m█[0m[38;2;133;199;201m█[0m[38;2;141;197;199m█[0m[38;2;140;197;199m█[0m");
$display("[38;2;219;209;130m█[0m[38;2;232;206;121m█[0m[38;2;240;208;107m█[0m[38;2;246;209;99m█[0m[38;2;254;214;94m█[0m[38;2;255;227;116m█[0m[38;2;252;228;122m█[0m[38;2;255;229;117m█[0m[38;2;253;225;120m█[0m[38;2;254;229;120m█[0m[38;2;255;227;119m█[0m[38;2;254;229;124m█[0m[38;2;253;229;124m█[0m[38;2;255;231;129m█[0m[38;2;254;217;95m█[0m[38;2;251;214;95m█[0m[38;2;247;214;109m█[0m[38;2;240;211;111m█[0m[38;2;224;208;120m█[0m[38;2;218;209;131m█[0m[38;2;209;209;136m█[0m[38;2;194;202;138m█[0m[38;2;182;202;151m█[0m[38;2;174;202;151m█[0m[38;2;170;197;154m█[0m[38;2;158;195;155m█[0m[38;2;158;197;165m█[0m[38;2;160;199;161m█[0m[38;2;161;198;156m█[0m[38;2;161;198;159m█[0m[38;2;161;201;161m█[0m[38;2;152;197;169m█[0m[38;2;150;197;165m█[0m[38;2;156;196;163m█[0m[38;2;138;192;164m█[0m[38;2;128;189;174m█[0m[38;2;121;192;183m█[0m[38;2;110;192;187m█[0m[38;2;106;186;185m█[0m[38;2;103;185;180m█[0m[38;2;96;188;188m█[0m[38;2;97;187;190m█[0m[38;2;95;187;189m█[0m[38;2;88;181;186m█[0m[38;2;89;184;192m█[0m[38;2;81;183;193m█[0m[38;2;76;181;193m█[0m[38;2;76;184;198m█[0m[38;2;66;178;195m█[0m[38;2;63;180;200m█[0m[38;2;55;178;199m█[0m[38;2;49;173;201m█[0m[38;2;42;174;200m█[0m[38;2;46;172;202m█[0m[38;2;43;171;199m█[0m[38;2;45;172;200m█[0m[38;2;45;172;201m█[0m[38;2;45;174;206m█[0m[38;2;40;170;203m█[0m[38;2;37;168;198m█[0m[38;2;41;172;203m█[0m[38;2;38;169;200m█[0m[38;2;36;169;199m█[0m[38;2;39;169;200m█[0m[38;2;37;167;198m█[0m[38;2;40;172;204m█[0m[38;2;42;175;206m█[0m[38;2;44;171;197m█[0m[38;2;115;202;210m█[0m[38;2;136;205;208m█[0m[38;2;169;216;208m█[0m[38;2;168;216;207m█[0m[38;2;189;218;207m█[0m[38;2;167;213;201m█[0m[38;2;184;221;208m█[0m[38;2;191;221;205m█[0m[38;2;177;218;209m█[0m[38;2;173;218;211m█[0m[38;2;156;217;209m█[0m[38;2;144;210;210m█[0m[38;2;140;209;209m█[0m[38;2;132;205;209m█[0m[38;2;126;206;212m█[0m[38;2;127;206;210m█[0m[38;2;121;204;210m█[0m[38;2;122;205;211m█[0m[38;2;122;206;210m█[0m[38;2;123;204;206m█[0m[38;2;135;206;210m█[0m[38;2;125;202;207m█[0m[38;2;129;203;205m█[0m[38;2;124;201;207m█[0m[38;2;126;201;206m█[0m[38;2;127;200;203m█[0m[38;2;126;198;206m█[0m[38;2;121;197;203m█[0m[38;2;122;195;202m█[0m[38;2;120;197;204m█[0m[38;2;113;194;207m█[0m[38;2;102;189;202m█[0m");
$display("[38;2;213;207;129m█[0m[38;2;223;205;124m█[0m[38;2;225;207;122m█[0m[38;2;224;207;122m█[0m[38;2;231;208;117m█[0m[38;2;244;212;107m█[0m[38;2;251;210;96m█[0m[38;2;252;210;94m█[0m[38;2;252;209;88m█[0m[38;2;253;211;86m█[0m[38;2;253;210;89m█[0m[38;2;253;213;91m█[0m[38;2;252;214;94m█[0m[38;2;243;210;105m█[0m[38;2;239;211;113m█[0m[38;2;225;207;119m█[0m[38;2;213;206;126m█[0m[38;2;217;207;128m█[0m[38;2;215;209;128m█[0m[38;2;215;206;127m█[0m[38;2;203;203;131m█[0m[38;2;187;203;145m█[0m[38;2;181;203;147m█[0m[38;2;177;204;153m█[0m[38;2;162;202;167m█[0m[38;2;140;194;171m█[0m[38;2;139;199;178m█[0m[38;2;129;195;175m█[0m[38;2;132;192;174m█[0m[38;2;130;196;179m█[0m[38;2;138;199;175m█[0m[38;2;143;195;170m█[0m[38;2;150;200;169m█[0m[38;2;145;196;170m█[0m[38;2;138;193;170m█[0m[38;2;132;193;173m█[0m[38;2;128;194;179m█[0m[38;2;115;189;178m█[0m[38;2;112;188;176m█[0m[38;2;126;196;180m█[0m[38;2;123;193;178m█[0m[38;2;112;190;180m█[0m[38;2;104;188;186m█[0m[38;2;105;190;188m█[0m[38;2;98;189;191m█[0m[38;2;91;188;192m█[0m[38;2;83;184;193m█[0m[38;2;81;186;196m█[0m[38;2;81;185;194m█[0m[38;2;80;184;195m█[0m[38;2;83;186;197m█[0m[38;2;77;185;200m█[0m[38;2;75;185;198m█[0m[38;2;78;185;196m█[0m[38;2;70;182;198m█[0m[38;2;63;182;203m█[0m[38;2;58;178;202m█[0m[38;2;55;179;203m█[0m[38;2;54;179;206m█[0m[38;2;47;174;201m█[0m[38;2;47;174;203m█[0m[38;2;46;176;203m█[0m[38;2;40;172;200m█[0m[38;2;39;171;200m█[0m[38;2;37;170;198m█[0m[38;2;39;170;201m█[0m[38;2;39;171;201m█[0m[38;2;41;172;200m█[0m[38;2;39;171;200m█[0m[38;2;43;173;208m█[0m[38;2;38;170;199m█[0m[38;2;42;176;203m█[0m[38;2;43;173;206m█[0m[38;2;49;178;202m█[0m[38;2;55;180;203m█[0m[38;2;46;171;205m█[0m[38;2;47;178;208m█[0m[38;2;55;178;205m█[0m[38;2;43;174;202m█[0m[38;2;45;173;200m█[0m[38;2;38;173;198m█[0m[38;2;44;172;205m█[0m[38;2;37;168;197m█[0m[38;2;41;170;199m█[0m[38;2;41;171;201m█[0m[38;2;39;166;202m█[0m[38;2;34;167;198m█[0m[38;2;39;174;206m█[0m[38;2;38;169;202m█[0m[38;2;37;169;201m█[0m[38;2;38;170;202m█[0m[38;2;36;164;198m█[0m[38;2;43;171;202m█[0m[38;2;41;170;200m█[0m[38;2;33;162;195m█[0m[38;2;39;172;203m█[0m[38;2;36;164;201m█[0m[38;2;36;166;199m█[0m[38;2;39;170;202m█[0m[38;2;41;171;201m█[0m");
$display("[38;2;207;207;138m█[0m[38;2;200;202;138m█[0m[38;2;199;205;138m█[0m[38;2;206;205;133m█[0m[38;2;212;204;129m█[0m[38;2;225;209;122m█[0m[38;2;228;211;122m█[0m[38;2;222;208;123m█[0m[38;2;211;204;127m█[0m[38;2;217;209;129m█[0m[38;2;230;208;119m█[0m[38;2;231;208;116m█[0m[38;2;228;209;120m█[0m[38;2;224;210;124m█[0m[38;2;218;209;129m█[0m[38;2;218;209;133m█[0m[38;2;205;205;137m█[0m[38;2;191;203;145m█[0m[38;2;186;202;147m█[0m[38;2;188;200;141m█[0m[38;2;189;203;143m█[0m[38;2;188;205;145m█[0m[38;2;187;203;147m█[0m[38;2;172;202;154m█[0m[38;2;160;199;160m█[0m[38;2;150;197;165m█[0m[38;2;145;197;171m█[0m[38;2;124;193;179m█[0m[38;2;108;192;188m█[0m[38;2;106;191;189m█[0m[38;2;103;192;192m█[0m[38;2;95;187;194m█[0m[38;2;97;191;188m█[0m[38;2;107;191;187m█[0m[38;2;107;191;186m█[0m[38;2;112;190;181m█[0m[38;2;122;191;176m█[0m[38;2;116;192;180m█[0m[38;2;120;194;185m█[0m[38;2;109;193;184m█[0m[38;2;103;189;186m█[0m[38;2;95;192;194m█[0m[38;2;90;190;195m█[0m[38;2;91;188;194m█[0m[38;2;89;189;193m█[0m[38;2;96;189;191m█[0m[38;2;108;194;189m█[0m[38;2;99;189;187m█[0m[38;2;92;187;190m█[0m[38;2;89;189;195m█[0m[38;2;90;189;199m█[0m[38;2;84;189;200m█[0m[38;2;80;185;194m█[0m[38;2;79;189;200m█[0m[38;2;71;185;198m█[0m[38;2;70;183;198m█[0m[38;2;71;187;203m█[0m[38;2;70;187;204m█[0m[38;2;69;183;199m█[0m[38;2;72;184;199m█[0m[38;2;66;182;199m█[0m[38;2;69;183;197m█[0m[38;2;56;178;199m█[0m[38;2;55;177;201m█[0m[38;2;53;177;201m█[0m[38;2;54;181;205m█[0m[38;2;53;179;204m█[0m[38;2;46;175;202m█[0m[38;2;47;177;201m█[0m[38;2;39;173;203m█[0m[38;2;45;176;206m█[0m[38;2;42;173;202m█[0m[38;2;39;172;203m█[0m[38;2;40;177;206m█[0m[38;2;39;170;201m█[0m[38;2;35;170;203m█[0m[38;2;37;172;201m█[0m[38;2;36;169;201m█[0m[38;2;41;174;207m█[0m[38;2;34;169;199m█[0m[38;2;37;171;202m█[0m[38;2;39;171;202m█[0m[38;2;37;169;200m█[0m[38;2;35;169;199m█[0m[38;2;31;166;198m█[0m[38;2;37;169;204m█[0m[38;2;33;166;201m█[0m[38;2;35;168;198m█[0m[38;2;33;168;200m█[0m[38;2;38;170;204m█[0m[38;2;34;168;199m█[0m[38;2;33;166;201m█[0m[38;2;34;166;199m█[0m[38;2;38;173;203m█[0m[38;2;35;168;202m█[0m[38;2;33;166;199m█[0m[38;2;31;166;196m█[0m[38;2;33;166;197m█[0m[38;2;34;166;197m█[0m[38;2;36;166;199m█[0m");
$display("[38;2;163;197;156m█[0m[38;2;171;200;149m█[0m[38;2;170;199;152m█[0m[38;2;186;203;146m█[0m[38;2;198;202;140m█[0m[38;2;211;207;131m█[0m[38;2;211;203;133m█[0m[38;2;196;203;138m█[0m[38;2;189;200;140m█[0m[38;2;190;201;138m█[0m[38;2;211;206;132m█[0m[38;2;206;203;130m█[0m[38;2;214;207;130m█[0m[38;2;222;209;129m█[0m[38;2;206;204;130m█[0m[38;2;194;201;138m█[0m[38;2;192;204;142m█[0m[38;2;179;201;143m█[0m[38;2;162;200;163m█[0m[38;2;150;197;168m█[0m[38;2;144;196;171m█[0m[38;2;171;202;160m█[0m[38;2;162;197;161m█[0m[38;2;171;200;155m█[0m[38;2;173;205;154m█[0m[38;2;165;199;155m█[0m[38;2;148;198;168m█[0m[38;2;139;199;176m█[0m[38;2;139;197;175m█[0m[38;2;129;194;178m█[0m[38;2;102;190;187m█[0m[38;2;94;189;192m█[0m[38;2;88;189;198m█[0m[38;2;83;190;198m█[0m[38;2;78;185;197m█[0m[38;2;85;191;198m█[0m[38;2;82;189;198m█[0m[38;2;85;189;196m█[0m[38;2;86;189;199m█[0m[38;2;87;190;195m█[0m[38;2;96;190;193m█[0m[38;2;104;194;192m█[0m[38;2;107;195;191m█[0m[38;2;100;195;196m█[0m[38;2;92;191;196m█[0m[38;2;90;193;201m█[0m[38;2;82;191;199m█[0m[38;2;82;191;204m█[0m[38;2;77;188;200m█[0m[38;2;83;188;201m█[0m[38;2;81;190;198m█[0m[38;2;94;187;192m█[0m[38;2;94;191;194m█[0m[38;2;98;192;194m█[0m[38;2;86;188;191m█[0m[38;2;83;189;195m█[0m[38;2;81;189;198m█[0m[38;2;75;188;200m█[0m[38;2;72;183;198m█[0m[38;2;74;188;204m█[0m[38;2;65;183;200m█[0m[38;2;72;189;208m█[0m[38;2;65;181;198m█[0m[38;2;62;182;202m█[0m[38;2;60;179;199m█[0m[38;2;58;179;202m█[0m[38;2;55;179;202m█[0m[38;2;58;188;206m█[0m[38;2;100;41;8m█[0m[38;2;85;39;8m█[0m[38;2;81;45;15m█[0m[38;2;80;44;7m█[0m[38;2;84;43;13m█[0m[38;2;50;178;193m█[0m[38;2;50;177;204m█[0m[38;2;44;170;199m█[0m[38;2;47;177;203m█[0m[38;2;43;177;207m█[0m[38;2;41;174;203m█[0m[38;2;41;176;202m█[0m[38;2;39;173;201m█[0m[38;2;38;171;201m█[0m[38;2;34;169;200m█[0m[38;2;29;165;197m█[0m[38;2;38;173;200m█[0m[38;2;37;168;199m█[0m[38;2;33;166;196m█[0m[38;2;33;167;199m█[0m[38;2;36;170;201m█[0m[38;2;32;166;196m█[0m[38;2;40;174;203m█[0m[38;2;32;166;197m█[0m[38;2;36;169;201m█[0m[38;2;35;166;201m█[0m[38;2;37;168;200m█[0m[38;2;37;170;202m█[0m[38;2;34;169;199m█[0m[38;2;32;168;201m█[0m[38;2;36;169;200m█[0m[38;2;37;169;197m█[0m");
$display("[38;2;138;198;172m█[0m[38;2;143;199;172m█[0m[38;2;160;197;162m█[0m[38;2;175;203;154m█[0m[38;2;190;205;147m█[0m[38;2;190;205;142m█[0m[38;2;193;205;145m█[0m[38;2;168;200;153m█[0m[38;2;163;196;157m█[0m[38;2;166;199;156m█[0m[38;2;169;204;159m█[0m[38;2;190;204;139m█[0m[38;2;188;204;147m█[0m[38;2;191;205;148m█[0m[38;2;205;206;134m█[0m[38;2;197;207;142m█[0m[38;2;176;202;152m█[0m[38;2;164;201;158m█[0m[38;2;161;202;158m█[0m[38;2;128;192;174m█[0m[38;2;125;196;179m█[0m[38;2;117;191;180m█[0m[38;2;124;198;184m█[0m[38;2;137;199;170m█[0m[38;2;139;199;173m█[0m[38;2;138;202;179m█[0m[38;2;142;198;174m█[0m[38;2;144;198;174m█[0m[38;2;135;201;184m█[0m[38;2;119;200;190m█[0m[38;2;108;194;190m█[0m[38;2;112;197;188m█[0m[38;2;113;198;192m█[0m[38;2;78;189;202m█[0m[38;2;76;192;205m█[0m[38;2;73;189;206m█[0m[38;2;66;189;201m█[0m[38;2;64;186;201m█[0m[38;2;67;190;205m█[0m[38;2;66;189;206m█[0m[38;2;71;188;203m█[0m[38;2;73;186;202m█[0m[38;2;73;189;202m█[0m[38;2;78;193;204m█[0m[38;2;88;196;203m█[0m[38;2;82;189;199m█[0m[38;2;84;190;197m█[0m[38;2;88;192;200m█[0m[38;2;87;195;204m█[0m[38;2;81;190;204m█[0m[38;2;77;190;199m█[0m[38;2;77;190;204m█[0m[38;2;74;189;203m█[0m[38;2;78;190;201m█[0m[38;2;70;184;200m█[0m[38;2;71;188;204m█[0m[38;2;75;186;202m█[0m[38;2;85;192;202m█[0m[38;2;77;189;200m█[0m[38;2;81;186;195m█[0m[38;2;76;186;198m█[0m[38;2;81;191;204m█[0m[38;2;71;184;199m█[0m[38;2;65;185;201m█[0m[38;2;97;107;95m█[0m[38;2;81;41;9m█[0m[38;2;89;48;13m█[0m[38;2;113;56;19m█[0m[38;2;252;213;125m█[0m[38;2;255;218;129m█[0m[38;2;254;221;134m█[0m[38;2;239;180;88m█[0m[38;2;75;38;12m█[0m[38;2;89;36;7m█[0m[38;2;56;176;197m█[0m[38;2;57;180;203m█[0m[38;2;49;175;198m█[0m[38;2;51;179;203m█[0m[38;2;47;177;205m█[0m[38;2;44;175;199m█[0m[38;2;40;173;199m█[0m[38;2;42;173;202m█[0m[38;2;44;177;206m█[0m[38;2;34;169;201m█[0m[38;2;37;171;200m█[0m[38;2;36;172;199m█[0m[38;2;37;171;200m█[0m[38;2;35;173;197m█[0m[38;2;41;176;204m█[0m[38;2;37;170;202m█[0m[38;2;39;173;199m█[0m[38;2;35;169;198m█[0m[38;2;42;171;201m█[0m[38;2;41;174;204m█[0m[38;2;37;169;197m█[0m[38;2;39;173;202m█[0m[38;2;42;173;201m█[0m[38;2;42;172;204m█[0m[38;2;40;172;199m█[0m[38;2;42;172;202m█[0m");
$display("[38;2;111;190;182m█[0m[38;2;129;197;182m█[0m[38;2;149;199;164m█[0m[38;2;156;198;161m█[0m[38;2;172;204;158m█[0m[38;2;159;195;154m█[0m[38;2;162;203;163m█[0m[38;2;142;196;169m█[0m[38;2;136;197;175m█[0m[38;2;141;195;169m█[0m[38;2;146;197;171m█[0m[38;2;172;200;156m█[0m[38;2;171;201;156m█[0m[38;2;177;204;155m█[0m[38;2;166;198;152m█[0m[38;2;178;203;149m█[0m[38;2;166;198;151m█[0m[38;2;146;199;172m█[0m[38;2;139;197;168m█[0m[38;2;138;197;168m█[0m[38;2;112;192;182m█[0m[38;2;103;191;188m█[0m[38;2;100;192;193m█[0m[38;2;96;192;192m█[0m[38;2;94;191;193m█[0m[38;2;116;197;188m█[0m[38;2;124;199;186m█[0m[38;2;119;197;188m█[0m[38;2;118;197;190m█[0m[38;2;122;198;183m█[0m[38;2;124;196;182m█[0m[38;2;97;195;194m█[0m[38;2;94;194;195m█[0m[38;2;97;197;198m█[0m[38;2;98;197;199m█[0m[38;2;85;194;201m█[0m[38;2;76;192;204m█[0m[38;2;70;191;205m█[0m[38;2;65;189;205m█[0m[38;2;67;191;208m█[0m[38;2;65;190;205m█[0m[38;2;63;192;207m█[0m[38;2;70;186;203m█[0m[38;2;68;191;203m█[0m[38;2;65;189;209m█[0m[38;2;68;185;207m█[0m[38;2;64;184;204m█[0m[38;2;66;189;206m█[0m[38;2;69;192;206m█[0m[38;2;73;189;198m█[0m[38;2;83;190;199m█[0m[38;2;81;190;204m█[0m[38;2;77;187;197m█[0m[38;2;78;189;204m█[0m[38;2;77;192;205m█[0m[38;2;67;187;201m█[0m[38;2;69;185;203m█[0m[38;2;71;190;204m█[0m[38;2;69;189;207m█[0m[38;2;69;187;207m█[0m[38;2;68;189;204m█[0m[38;2;76;189;206m█[0m[38;2;82;37;5m█[0m[38;2;88;44;12m█[0m[38;2;108;50;15m█[0m[38;2;255;216;124m█[0m[38;2;255;214;126m█[0m[38;2;226;168;75m█[0m[38;2;238;177;82m█[0m[38;2;243;183;91m█[0m[38;2;237;178;86m█[0m[38;2;241;180;89m█[0m[38;2;243;178;82m█[0m[38;2;81;42;11m█[0m[38;2;75;46;16m█[0m[38;2;52;177;203m█[0m[38;2;55;178;199m█[0m[38;2;51;175;199m█[0m[38;2;56;183;203m█[0m[38;2;48;179;201m█[0m[38;2;51;177;204m█[0m[38;2;46;175;205m█[0m[38;2;41;172;201m█[0m[38;2;42;175;203m█[0m[38;2;45;177;204m█[0m[38;2;43;175;205m█[0m[38;2;45;177;206m█[0m[38;2;45;176;203m█[0m[38;2;44;176;207m█[0m[38;2;44;174;202m█[0m[38;2;42;172;199m█[0m[38;2;39;171;199m█[0m[38;2;38;172;201m█[0m[38;2;45;174;201m█[0m[38;2;37;171;201m█[0m[38;2;45;177;202m█[0m[38;2;43;176;205m█[0m[38;2;45;174;200m█[0m[38;2;38;173;199m█[0m[38;2;48;175;204m█[0m");
$display("[38;2;96;194;193m█[0m[38;2;125;196;182m█[0m[38;2;133;198;174m█[0m[38;2;148;196;164m█[0m[38;2;148;199;169m█[0m[38;2;144;200;173m█[0m[38;2;133;196;175m█[0m[38;2;117;196;185m█[0m[38;2;117;196;187m█[0m[38;2;118;190;178m█[0m[38;2;126;195;176m█[0m[38;2;136;201;177m█[0m[38;2;160;201;164m█[0m[38;2;154;201;164m█[0m[38;2;153;198;164m█[0m[38;2;141;195;169m█[0m[38;2;153;197;157m█[0m[38;2;143;196;169m█[0m[38;2;121;192;177m█[0m[38;2;125;196;178m█[0m[38;2;120;196;183m█[0m[38;2;112;195;181m█[0m[38;2;92;192;194m█[0m[38;2;82;193;196m█[0m[38;2;80;191;200m█[0m[38;2;79;193;202m█[0m[38;2;79;189;197m█[0m[38;2;100;196;199m█[0m[38;2;109;197;193m█[0m[38;2;101;195;197m█[0m[38;2;101;198;200m█[0m[38;2;115;199;192m█[0m[38;2;114;197;192m█[0m[38;2;107;198;197m█[0m[38;2;93;194;197m█[0m[38;2;91;193;199m█[0m[38;2;96;200;203m█[0m[38;2;87;193;198m█[0m[38;2;71;190;204m█[0m[38;2;64;187;205m█[0m[38;2;65;189;206m█[0m[38;2;65;189;207m█[0m[38;2;63;190;209m█[0m[38;2;56;185;204m█[0m[38;2;65;189;211m█[0m[38;2;63;188;208m█[0m[38;2;63;188;206m█[0m[38;2;64;188;209m█[0m[38;2;61;188;206m█[0m[38;2;62;188;211m█[0m[38;2;68;190;208m█[0m[38;2;68;189;206m█[0m[38;2;71;185;199m█[0m[38;2;83;193;200m█[0m[38;2;84;191;199m█[0m[38;2;77;190;201m█[0m[38;2;76;190;201m█[0m[38;2;68;187;202m█[0m[38;2;68;186;207m█[0m[38;2;68;191;207m█[0m[38;2;92;46;11m█[0m[38;2;93;47;13m█[0m[38;2;255;230;137m█[0m[38;2;255;215;121m█[0m[38;2;254;212;121m█[0m[38;2;239;179;85m█[0m[38;2;242;181;86m█[0m[38;2;254;223;164m█[0m[38;2;255;243;215m█[0m[38;2;253;243;216m█[0m[38;2;244;182;86m█[0m[38;2;240;178;84m█[0m[38;2;237;177;83m█[0m[38;2;163;116;73m█[0m[38;2;77;39;12m█[0m[38;2;52;177;197m█[0m[38;2;51;176;205m█[0m[38;2;48;179;204m█[0m[38;2;41;175;202m█[0m[38;2;46;175;200m█[0m[38;2;48;179;204m█[0m[38;2;47;180;203m█[0m[38;2;46;176;204m█[0m[38;2;47;176;203m█[0m[38;2;41;174;200m█[0m[38;2;39;171;204m█[0m[38;2;43;173;200m█[0m[38;2;46;176;205m█[0m[38;2;47;180;207m█[0m[38;2;49;178;204m█[0m[38;2;43;176;205m█[0m[38;2;39;172;198m█[0m[38;2;43;175;204m█[0m[38;2;42;174;201m█[0m[38;2;45;175;205m█[0m[38;2;46;179;205m█[0m[38;2;50;179;201m█[0m[38;2;46;177;202m█[0m[38;2;45;177;202m█[0m[38;2;52;181;203m█[0m");
$display("[38;2;100;197;196m█[0m[38;2;113;197;188m█[0m[38;2;117;196;183m█[0m[38;2;170;216;203m█[0m[38;2;227;230;201m█[0m[38;2;227;231;201m█[0m[38;2;218;225;204m█[0m[38;2;188;218;199m█[0m[38;2;109;197;194m█[0m[38;2;114;197;191m█[0m[38;2;117;195;184m█[0m[38;2;114;197;185m█[0m[38;2;122;197;183m█[0m[38;2;139;200;177m█[0m[38;2;130;193;167m█[0m[38;2;132;198;177m█[0m[38;2;124;198;179m█[0m[38;2;141;199;170m█[0m[38;2;144;213;193m█[0m[38;2;107;195;187m█[0m[38;2;102;194;188m█[0m[38;2;101;194;192m█[0m[38;2;109;193;184m█[0m[38;2;88;198;203m█[0m[38;2;81;192;203m█[0m[38;2;76;192;205m█[0m[38;2;76;192;206m█[0m[38;2;68;193;204m█[0m[38;2;78;193;206m█[0m[38;2;87;194;202m█[0m[38;2;97;195;197m█[0m[38;2;89;198;206m█[0m[38;2;85;192;202m█[0m[38;2;99;198;203m█[0m[38;2;105;199;197m█[0m[38;2;106;199;195m█[0m[38;2;98;203;206m█[0m[38;2;91;195;202m█[0m[38;2;90;197;207m█[0m[38;2;84;191;200m█[0m[38;2;80;190;202m█[0m[38;2;64;191;210m█[0m[38;2;66;191;207m█[0m[38;2;64;189;205m█[0m[38;2;64;191;209m█[0m[38;2;60;186;209m█[0m[38;2;57;188;209m█[0m[38;2;58;187;205m█[0m[38;2;56;185;202m█[0m[38;2;55;185;205m█[0m[38;2;58;188;207m█[0m[38;2;68;189;212m█[0m[38;2;67;193;210m█[0m[38;2;68;191;209m█[0m[38;2;79;195;211m█[0m[38;2;72;187;201m█[0m[38;2;77;187;195m█[0m[38;2;77;194;202m█[0m[38;2;86;44;6m█[0m[38;2;87;43;11m█[0m[38;2;254;241;150m█[0m[38;2;255;210;117m█[0m[38;2;235;175;80m█[0m[38;2;245;186;89m█[0m[38;2;239;181;92m█[0m[38;2;254;245;220m█[0m[38;2;255;241;214m█[0m[38;2;254;242;217m█[0m[38;2;253;243;214m█[0m[38;2;255;242;218m█[0m[38;2;249;240;227m█[0m[38;2;240;179;85m█[0m[38;2;241;180;87m█[0m[38;2;235;175;93m█[0m[38;2;80;43;12m█[0m[38;2;42;21;11m█[0m[38;2;54;184;207m█[0m[38;2;54;183;204m█[0m[38;2;50;179;204m█[0m[38;2;50;181;204m█[0m[38;2;39;176;203m█[0m[38;2;43;178;206m█[0m[38;2;45;180;208m█[0m[38;2;48;182;204m█[0m[38;2;43;176;201m█[0m[38;2;39;175;204m█[0m[38;2;43;178;204m█[0m[38;2;40;178;201m█[0m[38;2;45;177;204m█[0m[38;2;41;176;201m█[0m[38;2;45;179;204m█[0m[38;2;47;182;206m█[0m[38;2;50;182;203m█[0m[38;2;47;179;201m█[0m[38;2;50;182;207m█[0m[38;2;45;178;203m█[0m[38;2;52;185;209m█[0m[38;2;46;182;203m█[0m[38;2;53;183;206m█[0m[38;2;57;184;204m█[0m");
$display("[38;2;96;195;197m█[0m[38;2;138;215;213m█[0m[38;2;194;224;205m█[0m[38;2;215;230;207m█[0m[38;2;221;231;206m█[0m[38;2;225;232;206m█[0m[38;2;228;232;205m█[0m[38;2;228;230;205m█[0m[38;2;226;233;205m█[0m[38;2;204;228;210m█[0m[38;2;103;194;189m█[0m[38;2;105;194;191m█[0m[38;2;106;196;191m█[0m[38;2;113;197;185m█[0m[38;2;121;195;180m█[0m[38;2;121;199;191m█[0m[38;2;117;197;183m█[0m[38;2;114;196;187m█[0m[38;2;133;198;175m█[0m[38;2;114;197;190m█[0m[38;2;100;196;194m█[0m[38;2;92;195;198m█[0m[38;2;99;193;194m█[0m[38;2;99;196;191m█[0m[38;2;77;191;200m█[0m[38;2;71;193;204m█[0m[38;2;71;194;209m█[0m[38;2;62;188;204m█[0m[38;2;64;190;209m█[0m[38;2;66;191;208m█[0m[38;2;69;196;209m█[0m[38;2;78;194;208m█[0m[38;2;88;196;203m█[0m[38;2;80;194;206m█[0m[38;2;83;192;201m█[0m[38;2;92;196;205m█[0m[38;2;96;195;198m█[0m[38;2;98;195;199m█[0m[38;2;93;196;198m█[0m[38;2;82;196;205m█[0m[38;2;77;194;206m█[0m[38;2;75;194;204m█[0m[38;2;81;195;208m█[0m[38;2;71;190;204m█[0m[38;2;62;189;207m█[0m[38;2;52;185;206m█[0m[38;2;53;188;209m█[0m[38;2;60;187;204m█[0m[38;2;54;187;209m█[0m[38;2;54;185;207m█[0m[38;2;51;183;206m█[0m[38;2;59;187;208m█[0m[38;2;59;191;210m█[0m[38;2;59;188;206m█[0m[38;2;43;80;70m█[0m[38;2;110;32;1m█[0m[38;2;90;42;5m█[0m[38;2;93;49;12m█[0m[38;2;92;46;11m█[0m[38;2;103;52;29m█[0m[38;2;69;20;0m█[0m[38;2;242;181;82m█[0m[38;2;236;181;88m█[0m[38;2;248;240;218m█[0m[38;2;255;242;217m█[0m[38;2;254;243;217m█[0m[38;2;254;241;215m█[0m[38;2;254;242;215m█[0m[38;2;253;241;216m█[0m[38;2;254;241;215m█[0m[38;2;255;242;210m█[0m[38;2;238;174;79m█[0m[38;2;237;176;83m█[0m[38;2;234;174;85m█[0m[38;2;71;37;16m█[0m[38;2;82;39;9m█[0m[38;2;68;189;205m█[0m[38;2;55;182;202m█[0m[38;2;57;185;205m█[0m[38;2;49;182;204m█[0m[38;2;51;183;206m█[0m[38;2;51;181;206m█[0m[38;2;47;181;204m█[0m[38;2;61;189;211m█[0m[38;2;49;182;207m█[0m[38;2;45;178;203m█[0m[38;2;48;183;207m█[0m[38;2;53;184;205m█[0m[38;2;51;182;208m█[0m[38;2;50;182;207m█[0m[38;2;51;183;207m█[0m[38;2;56;185;206m█[0m[38;2;53;183;202m█[0m[38;2;57;187;209m█[0m[38;2;60;186;205m█[0m[38;2;64;186;203m█[0m[38;2;61;186;204m█[0m[38;2;64;189;202m█[0m[38;2;65;191;207m█[0m[38;2;70;198;210m█[0m");
$display("[38;2;168;219;207m█[0m[38;2;174;223;209m█[0m[38;2;179;222;205m█[0m[38;2;185;225;207m█[0m[38;2;193;227;207m█[0m[38;2;180;225;212m█[0m[38;2;182;220;203m█[0m[38;2;195;228;212m█[0m[38;2;193;225;206m█[0m[38;2;196;225;206m█[0m[38;2;102;202;202m█[0m[38;2;92;194;195m█[0m[38;2;110;194;190m█[0m[38;2;104;199;196m█[0m[38;2;102;196;187m█[0m[38;2;103;196;188m█[0m[38;2;110;198;192m█[0m[38;2;102;196;190m█[0m[38;2;107;199;193m█[0m[38;2;127;197;177m█[0m[38;2;112;198;187m█[0m[38;2;92;191;192m█[0m[38;2;89;195;202m█[0m[38;2;93;195;195m█[0m[38;2;88;194;192m█[0m[38;2;73;192;205m█[0m[38;2;72;190;205m█[0m[38;2;65;191;207m█[0m[38;2;65;192;209m█[0m[38;2;60;191;209m█[0m[38;2;59;188;207m█[0m[38;2;63;191;207m█[0m[38;2;61;191;209m█[0m[38;2;70;192;200m█[0m[38;2;85;197;206m█[0m[38;2;78;196;208m█[0m[38;2;73;193;207m█[0m[38;2;88;198;201m█[0m[38;2;91;195;201m█[0m[38;2;100;198;201m█[0m[38;2;106;202;203m█[0m[38;2;85;194;201m█[0m[38;2;84;198;205m█[0m[38;2;79;195;205m█[0m[38;2;68;190;204m█[0m[38;2;70;193;210m█[0m[38;2;63;191;205m█[0m[38;2;67;189;207m█[0m[38;2;54;188;207m█[0m[38;2;115;46;10m█[0m[38;2;84;40;7m█[0m[38;2;90;45;14m█[0m[38;2;92;46;15m█[0m[38;2;95;50;14m█[0m[38;2;254;229;141m█[0m[38;2;253;197;84m█[0m[38;2;252;204;112m█[0m[38;2;253;203;109m█[0m[38;2;252;204;106m█[0m[38;2;255;204;108m█[0m[38;2;250;203;94m█[0m[38;2;254;198;89m█[0m[38;2;242;181;86m█[0m[38;2;239;176;83m█[0m[38;2;241;177;84m█[0m[38;2;226;164;73m█[0m[38;2;254;244;219m█[0m[38;2;254;242;214m█[0m[38;2;254;242;215m█[0m[38;2;255;241;215m█[0m[38;2;253;242;213m█[0m[38;2;242;182;85m█[0m[38;2;238;177;83m█[0m[38;2;236;174;81m█[0m[38;2;46;8;0m█[0m[38;2;77;39;13m█[0m[38;2;85;188;197m█[0m[38;2;66;185;198m█[0m[38;2;72;188;204m█[0m[38;2;64;189;206m█[0m[38;2;57;184;203m█[0m[38;2;56;182;205m█[0m[38;2;57;185;204m█[0m[38;2;54;182;205m█[0m[38;2;62;188;206m█[0m[38;2;59;185;206m█[0m[38;2;51;185;206m█[0m[38;2;56;185;205m█[0m[38;2;54;182;202m█[0m[38;2;57;183;203m█[0m[38;2;75;189;197m█[0m[38;2;65;188;201m█[0m[38;2;63;186;202m█[0m[38;2;67;190;204m█[0m[38;2;69;190;206m█[0m[38;2;67;189;202m█[0m[38;2;68;189;199m█[0m[38;2;67;187;199m█[0m[38;2;71;193;202m█[0m[38;2;76;196;205m█[0m");
$display("[38;2;166;221;208m█[0m[38;2;162;217;205m█[0m[38;2;149;217;211m█[0m[38;2;152;219;208m█[0m[38;2;154;216;209m█[0m[38;2;163;220;210m█[0m[38;2;160;218;209m█[0m[38;2;149;217;210m█[0m[38;2;156;219;212m█[0m[38;2;166;220;209m█[0m[38;2;156;215;208m█[0m[38;2;162;219;207m█[0m[38;2;177;226;212m█[0m[38;2;164;221;211m█[0m[38;2;153;217;207m█[0m[38;2;122;209;206m█[0m[38;2;128;211;208m█[0m[38;2;93;200;203m█[0m[38;2;85;194;196m█[0m[38;2;85;196;204m█[0m[38;2;103;38;2m█[0m[38;2;88;42;9m█[0m[38;2;91;48;10m█[0m[38;2;93;46;11m█[0m[38;2;93;45;12m█[0m[38;2;97;53;18m█[0m[38;2;75;23;4m█[0m[38;2;76;188;201m█[0m[38;2;74;195;206m█[0m[38;2;68;193;209m█[0m[38;2;61;191;211m█[0m[38;2;61;189;208m█[0m[38;2;62;189;207m█[0m[38;2;62;192;212m█[0m[38;2;53;185;200m█[0m[38;2;79;200;215m█[0m[38;2;77;199;210m█[0m[38;2;75;197;212m█[0m[38;2;74;194;210m█[0m[38;2;81;198;204m█[0m[38;2;93;197;197m█[0m[38;2;95;198;198m█[0m[38;2;89;198;203m█[0m[38;2;88;198;204m█[0m[38;2;80;191;202m█[0m[38;2;81;192;204m█[0m[38;2;83;40;7m█[0m[38;2;90;47;12m█[0m[38;2;97;51;11m█[0m[38;2;249;202;89m█[0m[38;2;255;205;102m█[0m[38;2;254;203;103m█[0m[38;2;254;204;101m█[0m[38;2;251;203;95m█[0m[38;2;237;178;83m█[0m[38;2;238;173;81m█[0m[38;2;238;179;84m█[0m[38;2;235;176;80m█[0m[38;2;239;175;85m█[0m[38;2;237;179;84m█[0m[38;2;233;174;79m█[0m[38;2;239;179;86m█[0m[38;2;236;174;80m█[0m[38;2;240;176;84m█[0m[38;2;238;180;85m█[0m[38;2;237;175;84m█[0m[38;2;239;177;84m█[0m[38;2;241;181;84m█[0m[38;2;236;176;80m█[0m[38;2;240;181;88m█[0m[38;2;240;180;85m█[0m[38;2;238;174;83m█[0m[38;2;240;180;85m█[0m[38;2;238;176;82m█[0m[38;2;244;199;130m█[0m[38;2;76;42;13m█[0m[38;2;94;185;194m█[0m[38;2;73;183;190m█[0m[38;2;78;192;201m█[0m[38;2;70;189;200m█[0m[38;2;71;187;199m█[0m[38;2;65;183;198m█[0m[38;2;71;190;204m█[0m[38;2;64;184;202m█[0m[38;2;59;186;204m█[0m[38;2;54;185;204m█[0m[38;2;61;187;206m█[0m[38;2;72;192;202m█[0m[38;2;66;187;204m█[0m[38;2;72;189;198m█[0m[38;2;79;191;195m█[0m[38;2;80;193;201m█[0m[38;2;86;189;195m█[0m[38;2;88;191;189m█[0m[38;2;85;190;186m█[0m[38;2;78;189;192m█[0m[38;2;80;190;191m█[0m[38;2;81;191;196m█[0m[38;2;88;190;194m█[0m[38;2;92;195;193m█[0m");
$display("[38;2;155;221;213m█[0m[38;2;147;217;212m█[0m[38;2;144;218;212m█[0m[38;2;142;214;209m█[0m[38;2;150;218;209m█[0m[38;2;142;213;208m█[0m[38;2;138;211;209m█[0m[38;2;136;216;209m█[0m[38;2;133;212;210m█[0m[38;2;128;208;206m█[0m[38;2;142;217;213m█[0m[38;2;128;210;212m█[0m[38;2;123;211;214m█[0m[38;2;115;210;212m█[0m[38;2;89;201;206m█[0m[38;2;93;196;207m█[0m[38;2;82;206;214m█[0m[38;2;94;46;11m█[0m[38;2;96;52;10m█[0m[38;2;99;45;12m█[0m[38;2;252;211;114m█[0m[38;2;255;215;117m█[0m[38;2;253;215;116m█[0m[38;2;253;204;100m█[0m[38;2;251;201;100m█[0m[38;2;253;207;105m█[0m[38;2;54;6;0m█[0m[38;2;90;46;12m█[0m[38;2;86;43;12m█[0m[38;2;70;182;194m█[0m[38;2;70;195;209m█[0m[38;2;62;191;209m█[0m[38;2;64;193;208m█[0m[38;2;61;191;208m█[0m[38;2;64;193;213m█[0m[38;2;64;193;214m█[0m[38;2;65;195;214m█[0m[38;2;70;195;212m█[0m[38;2;70;194;205m█[0m[38;2;64;191;207m█[0m[38;2;70;194;208m█[0m[38;2;72;194;208m█[0m[38;2;85;196;204m█[0m[38;2;95;197;208m█[0m[38;2;92;49;14m█[0m[38;2;93;50;10m█[0m[38;2;255;226;118m█[0m[38;2;254;205;104m█[0m[38;2;253;207;105m█[0m[38;2;252;205;100m█[0m[38;2;238;177;80m█[0m[38;2;240;175;85m█[0m[38;2;239;176;83m█[0m[38;2;238;174;81m█[0m[38;2;240;174;82m█[0m[38;2;239;178;86m█[0m[38;2;238;175;83m█[0m[38;2;241;181;87m█[0m[38;2;238;176;82m█[0m[38;2;241;180;88m█[0m[38;2;237;175;80m█[0m[38;2;238;177;85m█[0m[38;2;239;182;89m█[0m[38;2;241;177;86m█[0m[38;2;239;178;83m█[0m[38;2;237;175;83m█[0m[38;2;241;182;87m█[0m[38;2;242;183;90m█[0m[38;2;239;180;84m█[0m[38;2;240;181;87m█[0m[38;2;239;178;83m█[0m[38;2;238;180;84m█[0m[38;2;242;181;80m█[0m[38;2;78;37;6m█[0m[38;2;81;44;13m█[0m[38;2;75;38;8m█[0m[38;2;83;34;4m█[0m[38;2;85;184;196m█[0m[38;2;72;185;198m█[0m[38;2;72;189;201m█[0m[38;2;70;190;197m█[0m[38;2;70;190;201m█[0m[38;2;76;188;198m█[0m[38;2;71;188;204m█[0m[38;2;70;189;198m█[0m[38;2;66;191;206m█[0m[38;2;75;192;197m█[0m[38;2;66;186;200m█[0m[38;2;77;191;194m█[0m[38;2;77;190;200m█[0m[38;2;76;191;199m█[0m[38;2;83;190;192m█[0m[38;2;85;193;196m█[0m[38;2;98;196;187m█[0m[38;2;104;194;177m█[0m[38;2;104;199;182m█[0m[38;2;99;194;184m█[0m[38;2;110;196;176m█[0m[38;2;106;196;181m█[0m[38;2;115;201;177m█[0m");
$display("[38;2;80;193;205m█[0m[38;2;75;191;202m█[0m[38;2;90;193;197m█[0m[38;2;92;196;199m█[0m[38;2;92;197;197m█[0m[38;2;75;191;201m█[0m[38;2;72;189;203m█[0m[38;2;76;193;204m█[0m[38;2;73;190;202m█[0m[38;2;70;190;202m█[0m[38;2;67;191;206m█[0m[38;2;66;191;206m█[0m[38;2;73;189;199m█[0m[38;2;83;192;196m█[0m[38;2;62;194;208m█[0m[38;2;100;47;13m█[0m[38;2;106;54;12m█[0m[38;2;253;216;117m█[0m[38;2;255;216;120m█[0m[38;2;255;212;111m█[0m[38;2;238;176;84m█[0m[38;2;235;175;81m█[0m[38;2;243;181;90m█[0m[38;2;243;181;86m█[0m[38;2;241;182;89m█[0m[38;2;241;179;84m█[0m[38;2;240;179;83m█[0m[38;2;239;178;83m█[0m[38;2;72;29;7m█[0m[38;2;84;43;14m█[0m[38;2;88;200;205m█[0m[38;2;68;195;213m█[0m[38;2;67;194;211m█[0m[38;2;72;194;210m█[0m[38;2;72;199;213m█[0m[38;2;62;192;208m█[0m[38;2;69;195;211m█[0m[38;2;58;191;206m█[0m[38;2;60;192;213m█[0m[38;2;65;194;212m█[0m[38;2;73;195;211m█[0m[38;2;65;195;214m█[0m[38;2;82;45;10m█[0m[38;2;87;44;11m█[0m[38;2;254;238;142m█[0m[38;2;255;211;111m█[0m[38;2;253;210;107m█[0m[38;2;236;175;82m█[0m[38;2;240;180;88m█[0m[38;2;237;178;84m█[0m[38;2;237;176;80m█[0m[38;2;240;172;80m█[0m[38;2;236;177;84m█[0m[38;2;237;174;81m█[0m[38;2;238;175;81m█[0m[38;2;239;175;82m█[0m[38;2;238;177;83m█[0m[38;2;236;175;83m█[0m[38;2;238;178;84m█[0m[38;2;235;173;79m█[0m[38;2;240;178;87m█[0m[38;2;241;182;88m█[0m[38;2;239;178;82m█[0m[38;2;241;180;89m█[0m[38;2;239;174;81m█[0m[38;2;237;176;86m█[0m[38;2;239;176;82m█[0m[38;2;239;178;84m█[0m[38;2;239;178;80m█[0m[38;2;239;178;83m█[0m[38;2;241;179;87m█[0m[38;2;239;178;83m█[0m[38;2;237;175;82m█[0m[38;2;239;179;85m█[0m[38;2;237;178;85m█[0m[38;2;234;174;83m█[0m[38;2;252;208;116m█[0m[38;2;79;41;11m█[0m[38;2;79;41;14m█[0m[38;2;33;14;10m█[0m[38;2;71;188;197m█[0m[38;2;76;190;200m█[0m[38;2;73;188;203m█[0m[38;2;75;190;199m█[0m[38;2;83;193;195m█[0m[38;2;84;190;194m█[0m[38;2;88;193;188m█[0m[38;2;96;194;186m█[0m[38;2;99;197;186m█[0m[38;2;94;191;185m█[0m[38;2;88;191;190m█[0m[38;2;108;198;178m█[0m[38;2;111;197;176m█[0m[38;2;105;196;175m█[0m[38;2;110;198;178m█[0m[38;2;112;198;171m█[0m[38;2;113;200;173m█[0m[38;2;112;197;173m█[0m[38;2;118;198;171m█[0m[38;2;123;198;164m█[0m");
$display("[38;2;84;193;199m█[0m[38;2;90;193;198m█[0m[38;2;88;194;197m█[0m[38;2;83;188;190m█[0m[38;2;93;196;193m█[0m[38;2;81;191;198m█[0m[38;2;74;192;203m█[0m[38;2;72;190;200m█[0m[38;2;84;192;195m█[0m[38;2;79;194;201m█[0m[38;2;73;191;203m█[0m[38;2;75;193;200m█[0m[38;2;88;192;189m█[0m[38;2;56;23;7m█[0m[38;2;99;50;10m█[0m[38;2;255;238;141m█[0m[38;2;252;218;118m█[0m[38;2;241;180;86m█[0m[38;2;238;176;83m█[0m[38;2;239;177;83m█[0m[38;2;241;181;79m█[0m[38;2;205;148;81m█[0m[38;2;238;179;84m█[0m[38;2;240;179;83m█[0m[38;2;240;179;85m█[0m[38;2;235;170;79m█[0m[38;2;240;180;85m█[0m[38;2;238;178;85m█[0m[38;2;240;179;80m█[0m[38;2;89;43;8m█[0m[38;2;111;212;220m█[0m[38;2;67;192;212m█[0m[38;2;61;192;210m█[0m[38;2;67;195;211m█[0m[38;2;66;195;209m█[0m[38;2;71;198;215m█[0m[38;2;63;192;209m█[0m[38;2;59;191;209m█[0m[38;2;65;195;211m█[0m[38;2;67;199;218m█[0m[38;2;60;187;208m█[0m[38;2;84;41;8m█[0m[38;2;87;43;8m█[0m[38;2;255;212;110m█[0m[38;2;251;210;110m█[0m[38;2;236;175;81m█[0m[38;2;240;181;86m█[0m[38;2;245;179;87m█[0m[38;2;241;182;90m█[0m[38;2;238;179;85m█[0m[38;2;243;176;84m█[0m[38;2;230;181;76m█[0m[38;2;231;137;72m█[0m[38;2;249;175;94m█[0m[38;2;239;175;84m█[0m[38;2;237;178;85m█[0m[38;2;237;174;83m█[0m[38;2;238;174;80m█[0m[38;2;238;175;80m█[0m[38;2;237;176;82m█[0m[38;2;236;176;85m█[0m[38;2;238;176;79m█[0m[38;2;238;176;82m█[0m[38;2;239;179;85m█[0m[38;2;235;174;79m█[0m[38;2;236;175;84m█[0m[38;2;237;179;86m█[0m[38;2;240;177;85m█[0m[38;2;236;177;82m█[0m[38;2;239;176;85m█[0m[38;2;241;179;79m█[0m[38;2;74;35;6m█[0m[38;2;255;212;121m█[0m[38;2;240;176;85m█[0m[38;2;237;176;82m█[0m[38;2;240;181;86m█[0m[38;2;238;180;86m█[0m[38;2;239;181;87m█[0m[38;2;239;177;85m█[0m[38;2;77;43;15m█[0m[38;2;74;39;10m█[0m[38;2;56;5;0m█[0m[38;2;76;188;200m█[0m[38;2;73;184;189m█[0m[38;2;84;191;198m█[0m[38;2;93;194;192m█[0m[38;2;93;194;184m█[0m[38;2;92;191;185m█[0m[38;2;89;192;186m█[0m[38;2;99;195;188m█[0m[38;2;99;192;174m█[0m[38;2;103;195;176m█[0m[38;2;113;197;173m█[0m[38;2;109;197;168m█[0m[38;2;114;200;175m█[0m[38;2;114;197;166m█[0m[38;2;116;197;164m█[0m[38;2;112;195;164m█[0m[38;2;113;194;161m█[0m[38;2;120;200;167m█[0m");
$display("[38;2;109;201;189m█[0m[38;2;96;194;186m█[0m[38;2;103;194;180m█[0m[38;2;99;194;181m█[0m[38;2;104;198;189m█[0m[38;2;90;193;192m█[0m[38;2;91;192;192m█[0m[38;2;100;198;185m█[0m[38;2;94;191;188m█[0m[38;2;88;193;194m█[0m[38;2;89;194;195m█[0m[38;2;107;200;183m█[0m[38;2;106;223;221m█[0m[38;2;93;47;10m█[0m[38;2;246;202;104m█[0m[38;2;238;186;88m█[0m[38;2;238;178;82m█[0m[38;2;237;178;83m█[0m[38;2;227;175;90m█[0m[38;2;93;45;10m█[0m[38;2;100;52;26m█[0m[38;2;240;177;84m█[0m[38;2;241;180;88m█[0m[38;2;242;181;88m█[0m[38;2;255;217;130m█[0m[38;2;92;50;21m█[0m[38;2;89;44;7m█[0m[38;2;87;43;13m█[0m[38;2;89;45;13m█[0m[38;2;89;46;14m█[0m[38;2;88;45;12m█[0m[38;2;91;46;14m█[0m[38;2;86;47;12m█[0m[38;2;95;46;16m█[0m[38;2;87;43;13m█[0m[38;2;88;43;11m█[0m[38;2;77;47;14m█[0m[38;2;92;34;1m█[0m[38;2;109;159;158m█[0m[38;2;70;189;204m█[0m[38;2;75;35;7m█[0m[38;2;90;45;7m█[0m[38;2;255;208;108m█[0m[38;2;236;169;69m█[0m[38;2;255;242;207m█[0m[38;2;254;238;208m█[0m[38;2;253;237;207m█[0m[38;2;252;238;206m█[0m[38;2;253;237;205m█[0m[38;2;253;236;207m█[0m[38;2;240;134;94m█[0m[38;2;241;138;98m█[0m[38;2;241;136;96m█[0m[38;2;239;135;92m█[0m[38;2;242;129;89m█[0m[38;2;244;130;88m█[0m[38;2;234;131;78m█[0m[38;2;242;176;83m█[0m[38;2;240;180;87m█[0m[38;2;239;180;88m█[0m[38;2;238;177;85m█[0m[38;2;237;173;90m█[0m[38;2;242;181;87m█[0m[38;2;242;183;89m█[0m[38;2;244;180;87m█[0m[38;2;239;179;85m█[0m[38;2;237;175;82m█[0m[38;2;240;176;81m█[0m[38;2;240;179;85m█[0m[38;2;239;181;88m█[0m[38;2;240;181;88m█[0m[38;2;50;16;3m█[0m[38;2;81;44;11m█[0m[38;2;234;177;79m█[0m[38;2;239;176;84m█[0m[38;2;238;178;84m█[0m[38;2;238;181;89m█[0m[38;2;239;180;85m█[0m[38;2;240;177;83m█[0m[38;2;239;181;84m█[0m[38;2;241;180;84m█[0m[38;2;76;41;14m█[0m[38;2;67;38;12m█[0m[38;2;82;188;191m█[0m[38;2;89;195;186m█[0m[38;2;95;192;187m█[0m[38;2;98;192;178m█[0m[38;2;102;195;177m█[0m[38;2;103;194;176m█[0m[38;2;104;194;174m█[0m[38;2;110;196;173m█[0m[38;2;104;192;171m█[0m[38;2;112;197;164m█[0m[38;2;111;197;164m█[0m[38;2;113;192;162m█[0m[38;2;113;196;160m█[0m[38;2;117;196;161m█[0m[38;2;114;199;168m█[0m[38;2;111;194;161m█[0m[38;2;122;199;157m█[0m");
$display("[38;2;114;196;169m█[0m[38;2;113;192;167m█[0m[38;2;113;197;170m█[0m[38;2;116;197;168m█[0m[38;2;112;197;171m█[0m[38;2;104;195;168m█[0m[38;2;114;198;168m█[0m[38;2;116;200;173m█[0m[38;2;111;202;181m█[0m[38;2;102;196;185m█[0m[38;2;113;196;176m█[0m[38;2;125;198;172m█[0m[38;2;96;43;11m█[0m[38;2;62;22;0m█[0m[38;2;244;181;86m█[0m[38;2;236;177;81m█[0m[38;2;239;181;88m█[0m[38;2;245;189;96m█[0m[38;2;96;51;13m█[0m[38;2;255;215;120m█[0m[38;2;166;111;43m█[0m[38;2;90;44;12m█[0m[38;2;92;46;13m█[0m[38;2;95;48;10m█[0m[38;2;130;71;21m█[0m[38;2;254;208;112m█[0m[38;2;255;203;103m█[0m[38;2;254;205;104m█[0m[38;2;254;203;100m█[0m[38;2;251;199;97m█[0m[38;2;253;202;99m█[0m[38;2;252;201;98m█[0m[38;2;255;203;98m█[0m[38;2;253;200;97m█[0m[38;2;238;174;76m█[0m[38;2;241;179;87m█[0m[38;2;239;172;76m█[0m[38;2;243;178;87m█[0m[38;2;176;119;65m█[0m[38;2;83;40;10m█[0m[38;2;84;42;12m█[0m[38;2;77;28;0m█[0m[38;2;254;237;207m█[0m[38;2;254;238;207m█[0m[38;2;255;241;210m█[0m[38;2;255;236;208m█[0m[38;2;255;241;208m█[0m[38;2;253;238;208m█[0m[38;2;253;239;206m█[0m[38;2;250;236;204m█[0m[38;2;239;132;97m█[0m[38;2;245;135;97m█[0m[38;2;239;132;91m█[0m[38;2;244;137;98m█[0m[38;2;244;137;97m█[0m[38;2;250;242;209m█[0m[38;2;243;137;91m█[0m[38;2;246;129;92m█[0m[38;2;237;176;82m█[0m[38;2;237;173;82m█[0m[38;2;255;216;129m█[0m[38;2;79;37;7m█[0m[38;2;71;36;16m█[0m[38;2;240;177;85m█[0m[38;2;236;173;84m█[0m[38;2;238;178;86m█[0m[38;2;239;174;80m█[0m[38;2;233;173;78m█[0m[38;2;238;177;84m█[0m[38;2;240;180;87m█[0m[38;2;240;177;86m█[0m[38;2;242;180;89m█[0m[38;2;236;176;85m█[0m[38;2;235;174;78m█[0m[38;2;239;181;87m█[0m[38;2;237;179;84m█[0m[38;2;238;179;87m█[0m[38;2;239;179;83m█[0m[38;2;236;177;83m█[0m[38;2;241;180;85m█[0m[38;2;240;181;86m█[0m[38;2;239;184;88m█[0m[38;2;79;39;9m█[0m[38;2;75;37;8m█[0m[38;2;75;38;13m█[0m[38;2;76;41;14m█[0m[38;2;77;41;9m█[0m[38;2;75;44;9m█[0m[38;2;96;38;18m█[0m[38;2;155;231;199m█[0m[38;2;114;192;158m█[0m[38;2;115;195;157m█[0m[38;2;114;196;156m█[0m[38;2;115;196;158m█[0m[38;2;115;195;158m█[0m[38;2;116;195;158m█[0m[38;2;107;192;157m█[0m[38;2;116;195;159m█[0m[38;2;114;194;151m█[0m[38;2;109;193;154m█[0m");
$display("[38;2;122;196;155m█[0m[38;2;119;193;155m█[0m[38;2;121;193;155m█[0m[38;2;112;192;157m█[0m[38;2;115;192;153m█[0m[38;2;120;198;162m█[0m[38;2;124;195;155m█[0m[38;2;120;195;153m█[0m[38;2;127;198;157m█[0m[38;2;121;197;160m█[0m[38;2;123;198;157m█[0m[38;2;156;223;183m█[0m[38;2;86;42;14m█[0m[38;2;244;184;83m█[0m[38;2;239;181;86m█[0m[38;2;240;180;86m█[0m[38;2;237;174;81m█[0m[38;2;255;202;102m█[0m[38;2;90;44;8m█[0m[38;2;97;48;16m█[0m[38;2;90;35;7m█[0m[38;2;255;210;112m█[0m[38;2;255;207;108m█[0m[38;2;252;205;101m█[0m[38;2;252;203;100m█[0m[38;2;241;182;89m█[0m[38;2;237;178;82m█[0m[38;2;237;174;82m█[0m[38;2;239;180;87m█[0m[38;2;239;177;82m█[0m[38;2;240;176;85m█[0m[38;2;240;172;81m█[0m[38;2;240;177;77m█[0m[38;2;84;43;14m█[0m[38;2;84;44;11m█[0m[38;2;82;41;12m█[0m[38;2;83;44;13m█[0m[38;2;47;13;0m█[0m[38;2;239;180;88m█[0m[38;2;255;210;119m█[0m[38;2;85;42;10m█[0m[38;2;252;236;205m█[0m[38;2;253;236;205m█[0m[38;2;252;237;206m█[0m[38;2;255;239;210m█[0m[38;2;254;236;205m█[0m[38;2;254;238;207m█[0m[38;2;255;238;207m█[0m[38;2;254;239;208m█[0m[38;2;254;238;206m█[0m[38;2;254;240;210m█[0m[38;2;247;236;221m█[0m[38;2;239;142;98m█[0m[38;2;241;134;94m█[0m[38;2;241;135;94m█[0m[38;2;244;131;90m█[0m[38;2;240;129;88m█[0m[38;2;234;128;87m█[0m[38;2;240;178;79m█[0m[38;2;234;171;79m█[0m[38;2;239;177;84m█[0m[38;2;235;174;80m█[0m[38;2;46;5;0m█[0m[38;2;82;43;16m█[0m[38;2;84;45;14m█[0m[38;2;79;40;9m█[0m[38;2;237;178;87m█[0m[38;2;238;175;81m█[0m[38;2;235;178;81m█[0m[38;2;240;180;87m█[0m[38;2;238;177;82m█[0m[38;2;237;175;81m█[0m[38;2;239;179;83m█[0m[38;2;239;176;81m█[0m[38;2;234;176;82m█[0m[38;2;241;181;83m█[0m[38;2;240;179;85m█[0m[38;2;235;177;81m█[0m[38;2;236;173;79m█[0m[38;2;239;178;85m█[0m[38;2;238;176;84m█[0m[38;2;242;182;89m█[0m[38;2;236;174;67m█[0m[38;2;80;40;4m█[0m[38;2;233;174;78m█[0m[38;2;235;173;81m█[0m[38;2;234;175;82m█[0m[38;2;237;177;85m█[0m[38;2;242;180;88m█[0m[38;2;165;111;32m█[0m[38;2;75;40;10m█[0m[38;2;75;35;5m█[0m[38;2;76;40;13m█[0m[38;2;75;39;10m█[0m[38;2;103;206;151m█[0m[38;2;116;192;146m█[0m[38;2;110;190;148m█[0m[38;2;107;189;151m█[0m[38;2;109;188;147m█[0m[38;2;108;187;149m█[0m");
$display("[38;2;134;197;139m█[0m[38;2;123;191;146m█[0m[38;2;121;191;143m█[0m[38;2;132;196;139m█[0m[38;2;130;195;142m█[0m[38;2;123;192;140m█[0m[38;2;126;196;148m█[0m[38;2;127;197;151m█[0m[38;2;135;200;141m█[0m[38;2;136;199;144m█[0m[38;2;131;194;138m█[0m[38;2;171;223;176m█[0m[38;2;85;41;10m█[0m[38;2;218;148;50m█[0m[38;2;235;175;80m█[0m[38;2;239;176;80m█[0m[38;2;90;45;7m█[0m[38;2;97;51;14m█[0m[38;2;254;238;135m█[0m[38;2;253;209;109m█[0m[38;2;250;207;107m█[0m[38;2;238;177;84m█[0m[38;2;240;177;84m█[0m[38;2;242;180;86m█[0m[38;2;240;175;85m█[0m[38;2;236;175;80m█[0m[38;2;238;177;84m█[0m[38;2;235;173;79m█[0m[38;2;238;178;84m█[0m[38;2;236;176;80m█[0m[38;2;237;175;85m█[0m[38;2;82;41;11m█[0m[38;2;85;43;9m█[0m[38;2;247;238;209m█[0m[38;2;254;240;209m█[0m[38;2;255;239;209m█[0m[38;2;254;237;205m█[0m[38;2;97;51;13m█[0m[38;2;86;43;13m█[0m[38;2;80;39;10m█[0m[38;2;87;44;13m█[0m[38;2;255;239;208m█[0m[38;2;255;239;206m█[0m[38;2;254;237;206m█[0m[38;2;254;238;208m█[0m[38;2;253;237;208m█[0m[38;2;254;238;207m█[0m[38;2;253;241;209m█[0m[38;2;254;239;207m█[0m[38;2;253;237;207m█[0m[38;2;254;238;208m█[0m[38;2;255;238;208m█[0m[38;2;252;238;206m█[0m[38;2;252;235;204m█[0m[38;2;252;239;207m█[0m[38;2;248;236;208m█[0m[38;2;255;237;208m█[0m[38;2;253;234;204m█[0m[38;2;254;238;207m█[0m[38;2;221;162;70m█[0m[38;2;234;178;88m█[0m[38;2;235;173;79m█[0m[38;2;236;177;85m█[0m[38;2;237;178;85m█[0m[38;2;232;173;80m█[0m[38;2;237;176;81m█[0m[38;2;236;176;81m█[0m[38;2;237;176;82m█[0m[38;2;236;176;83m█[0m[38;2;233;170;77m█[0m[38;2;237;176;83m█[0m[38;2;235;173;82m█[0m[38;2;242;180;86m█[0m[38;2;234;178;82m█[0m[38;2;241;180;84m█[0m[38;2;235;175;79m█[0m[38;2;239;179;85m█[0m[38;2;73;41;12m█[0m[38;2;79;42;9m█[0m[38;2;237;175;83m█[0m[38;2;240;178;84m█[0m[38;2;237;176;81m█[0m[38;2;235;176;79m█[0m[38;2;236;172;78m█[0m[38;2;238;178;84m█[0m[38;2;221;173;105m█[0m[38;2;216;162;71m█[0m[38;2;243;174;77m█[0m[38;2;241;177;80m█[0m[38;2;234;178;83m█[0m[38;2;235;174;81m█[0m[38;2;236;177;81m█[0m[38;2;239;178;87m█[0m[38;2;243;182;90m█[0m[38;2;75;41;14m█[0m[38;2;83;39;13m█[0m[38;2;120;187;139m█[0m[38;2;104;184;141m█[0m[38;2;103;185;139m█[0m[38;2;108;185;138m█[0m");
$display("[38;2;112;180;130m█[0m[38;2;106;175;127m█[0m[38;2;114;179;126m█[0m[38;2;107;176;128m█[0m[38;2;120;189;135m█[0m[38;2;122;189;137m█[0m[38;2;127;192;136m█[0m[38;2;134;192;131m█[0m[38;2;137;198;134m█[0m[38;2;128;193;135m█[0m[38;2;126;190;129m█[0m[38;2;120;189;134m█[0m[38;2;83;37;11m█[0m[38;2;62;26;10m█[0m[38;2;227;164;84m█[0m[38;2;90;43;12m█[0m[38;2;63;18;0m█[0m[38;2;255;207;105m█[0m[38;2;255;216;120m█[0m[38;2;238;176;83m██[0m[38;2;242;180;87m█[0m[38;2;239;177;86m█[0m[38;2;240;180;86m█[0m[38;2;236;176;82m█[0m[38;2;238;178;82m█[0m[38;2;240;176;85m█[0m[38;2;238;175;81m█[0m[38;2;239;176;83m█[0m[38;2;236;172;80m█[0m[38;2;87;46;13m█[0m[38;2;89;40;11m█[0m[38;2;255;240;210m█[0m[38;2;255;239;210m█[0m[38;2;255;240;210m█[0m[38;2;254;240;209m█[0m[38;2;253;236;205m█[0m[38;2;254;239;208m█[0m[38;2;253;236;207m█[0m[38;2;90;48;16m█[0m[38;2;89;45;16m█[0m[38;2;252;239;209m█[0m[38;2;254;239;209m█[0m[38;2;255;239;208m█[0m[38;2;255;238;208m█[0m[38;2;255;240;208m█[0m[38;2;254;236;206m█[0m[38;2;254;235;206m█[0m[38;2;252;237;203m█[0m[38;2;254;236;206m█[0m[38;2;254;239;208m█[0m[38;2;255;240;208m█[0m[38;2;255;239;206m█[0m[38;2;254;236;204m█[0m[38;2;252;234;205m█[0m[38;2;253;237;206m█[0m[38;2;254;240;209m█[0m[38;2;254;238;205m█[0m[38;2;254;237;205m█[0m[38;2;255;238;210m█[0m[38;2;254;235;206m█[0m[38;2;253;235;211m█[0m[38;2;255;241;190m█[0m[38;2;243;177;76m█[0m[38;2;235;174;79m█[0m[38;2;237;174;79m█[0m[38;2;236;171;80m█[0m[38;2;233;172;78m█[0m[38;2;236;173;77m█[0m[38;2;235;173;78m█[0m[38;2;233;174;81m█[0m[38;2;235;174;80m█[0m[38;2;241;180;85m█[0m[38;2;236;176;83m█[0m[38;2;237;177;86m█[0m[38;2;239;179;86m█[0m[38;2;241;179;84m█[0m[38;2;235;175;89m█[0m[38;2;73;35;4m█[0m[38;2;236;177;83m█[0m[38;2;236;179;84m█[0m[38;2;239;179;84m█[0m[38;2;242;182;87m█[0m[38;2;236;177;81m█[0m[38;2;241;173;77m█[0m[38;2;253;240;210m█[0m[38;2;254;239;210m█[0m[38;2;253;241;211m█[0m[38;2;254;238;212m█[0m[38;2;255;240;208m█[0m[38;2;255;242;215m█[0m[38;2;214;161;76m█[0m[38;2;233;173;79m█[0m[38;2;238;180;85m█[0m[38;2;73;38;16m█[0m[38;2;73;36;11m█[0m[38;2;96;176;134m█[0m[38;2;100;180;132m█[0m[38;2;91;175;128m█[0m[38;2;96;178;130m█[0m");
$display("[38;2;95;168;120m█[0m[38;2;90;167;121m█[0m[38;2;92;165;116m█[0m[38;2;92;166;116m█[0m[38;2;91;165;115m█[0m[38;2;100;171;113m█[0m[38;2;122;185;120m█[0m[38;2;101;171;119m█[0m[38;2;94;168;122m█[0m[38;2;103;175;123m█[0m[38;2;101;171;117m█[0m[38;2;113;181;122m█[0m[38;2;142;228;167m█[0m[38;2;77;39;12m█[0m[38;2;96;50;14m█[0m[38;2;249;204;93m█[0m[38;2;254;211;112m█[0m[38;2;245;183;90m█[0m[38;2;241;180;83m█[0m[38;2;238;179;84m█[0m[38;2;237;175;81m█[0m[38;2;236;172;78m█[0m[38;2;241;181;87m█[0m[38;2;238;176;80m█[0m[38;2;237;174;79m█[0m[38;2;237;179;86m█[0m[38;2;237;176;82m█[0m[38;2;238;175;83m█[0m[38;2;239;176;84m█[0m[38;2;239;174;84m█[0m[38;2;83;42;11m█[0m[38;2;32;0;0m█[0m[38;2;252;238;207m█[0m[38;2;254;237;206m█[0m[38;2;254;238;207m█[0m[38;2;254;238;206m█[0m[38;2;255;239;210m█[0m[38;2;254;237;206m█[0m[38;2;252;237;206m█[0m[38;2;251;253;238m█[0m[38;2;88;44;14m█[0m[38;2;252;255;244m█[0m[38;2;254;238;208m█[0m[38;2;253;237;208m█[0m[38;2;255;237;205m█[0m[38;2;253;238;208m█[0m[38;2;254;236;205m█[0m[38;2;254;236;208m█[0m[38;2;255;240;210m█[0m[38;2;255;237;209m█[0m[38;2;254;237;204m█[0m[38;2;253;239;208m█[0m[38;2;253;238;209m█[0m[38;2;252;237;207m█[0m[38;2;255;239;206m█[0m[38;2;254;238;205m█[0m[38;2;253;235;207m█[0m[38;2;254;237;207m█[0m[38;2;252;235;205m█[0m[38;2;254;238;204m█[0m[38;2;253;236;204m█[0m[38;2;254;236;207m█[0m[38;2;254;237;204m█[0m[38;2;252;237;205m█[0m[38;2;254;238;206m█[0m[38;2;249;255;247m█[0m[38;2;80;44;13m█[0m[38;2;84;45;22m█[0m[38;2;76;39;11m█[0m[38;2;80;40;12m█[0m[38;2;238;175;82m█[0m[38;2;242;181;88m█[0m[38;2;237;176;83m█[0m[38;2;237;178;83m█[0m[38;2;236;177;83m█[0m[38;2;239;177;84m█[0m[38;2;245;186;88m█[0m[38;2;239;179;85m█[0m[38;2;236;176;82m█[0m[38;2;237;176;81m█[0m[38;2;239;175;84m█[0m[38;2;238;177;84m█[0m[38;2;238;177;85m█[0m[38;2;239;176;84m█[0m[38;2;237;176;85m█[0m[38;2;248;236;219m█[0m[38;2;254;238;210m█[0m[38;2;255;240;209m██[0m[38;2;255;240;213m█[0m[38;2;254;240;215m█[0m[38;2;238;173;81m█[0m[38;2;233;171;80m█[0m[38;2;73;29;0m█[0m[38;2;73;37;9m█[0m[38;2;94;180;132m█[0m[38;2;81;168;122m█[0m[38;2;82;164;117m█[0m[38;2;80;164;111m█[0m[38;2;73;159;116m█[0m");
$display("[38;2;86;161;110m█[0m[38;2;84;162;110m█[0m[38;2;84;158;109m█[0m[38;2;88;165;115m█[0m[38;2;89;162;108m█[0m[38;2;92;170;120m█[0m[38;2;79;159;114m█[0m[38;2;90;167;116m█[0m[38;2;86;164;113m█[0m[38;2;79;158;107m█[0m[38;2;83;162;114m█[0m[38;2;77;157;106m█[0m[38;2;47;28;0m█[0m[38;2;88;45;12m█[0m[38;2;249;208;100m█[0m[38;2;254;213;109m█[0m[38;2;242;180;85m█[0m[38;2;243;183;88m█[0m[38;2;236;176;78m█[0m[38;2;240;179;85m█[0m[38;2;238;176;84m█[0m[38;2;236;175;83m█[0m[38;2;239;175;83m█[0m[38;2;235;174;78m█[0m[38;2;239;176;82m█[0m[38;2;236;177;82m█[0m[38;2;237;176;82m█[0m[38;2;235;175;78m█[0m[38;2;239;178;84m█[0m[38;2;240;179;85m█[0m[38;2;68;30;4m█[0m[38;2;84;43;15m█[0m[38;2;248;234;206m█[0m[38;2;255;240;210m█[0m[38;2;254;240;210m█[0m[38;2;254;237;206m█[0m[38;2;254;238;206m█[0m[38;2;253;238;206m█[0m[38;2;255;238;210m█[0m[38;2;254;237;204m█[0m[38;2;86;42;14m█[0m[38;2;75;34;12m█[0m[38;2;255;239;211m█[0m[38;2;254;240;209m█[0m[38;2;255;240;211m█[0m[38;2;253;239;209m█[0m[38;2;255;237;209m█[0m[38;2;253;238;208m█[0m[38;2;252;239;206m█[0m[38;2;254;237;206m█[0m[38;2;255;238;207m█[0m[38;2;254;239;206m█[0m[38;2;254;236;206m█[0m[38;2;254;237;207m█[0m[38;2;253;238;206m█[0m[38;2;254;237;208m█[0m[38;2;255;239;207m█[0m[38;2;250;234;205m█[0m[38;2;250;235;204m█[0m[38;2;73;38;11m█[0m[38;2;253;248;233m█[0m[38;2;255;234;205m█[0m[38;2;254;238;204m█[0m[38;2;254;236;206m█[0m[38;2;255;237;207m█[0m[38;2;253;239;207m█[0m[38;2;77;39;12m█[0m[38;2;74;38;10m█[0m[38;2;75;39;11m█[0m[38;2;74;35;11m█[0m[38;2;69;34;5m█[0m[38;2;237;180;90m█[0m[38;2;240;183;89m█[0m[38;2;236;179;84m█[0m[38;2;236;176;80m█[0m[38;2;240;180;88m█[0m[38;2;239;178;86m█[0m[38;2;238;179;85m█[0m[38;2;235;175;79m█[0m[38;2;241;181;86m█[0m[38;2;240;179;86m█[0m[38;2;240;178;84m█[0m[38;2;240;180;86m█[0m[38;2;235;174;82m█[0m[38;2;232;172;78m█[0m[38;2;234;173;78m█[0m[38;2;254;240;212m█[0m[38;2;254;239;210m█[0m[38;2;254;238;211m█[0m[38;2;241;174;71m█[0m[38;2;235;174;79m█[0m[38;2;234;175;85m█[0m[38;2;60;28;8m█[0m[38;2;73;36;10m█[0m[38;2;69;175;132m█[0m[38;2;69;157;114m█[0m[38;2;71;155;107m█[0m[38;2;62;151;105m█[0m[38;2;69;152;104m█[0m[38;2;58;148;105m█[0m");
$display("[38;2;88;161;102m█[0m[38;2;90;162;99m█[0m[38;2;119;182;94m█[0m[38;2;109;170;87m█[0m[38;2;93;167;99m█[0m[38;2;118;172;65m█[0m[38;2;76;157;105m█[0m[38;2;84;160;102m█[0m[38;2;81;159;97m█[0m[38;2;85;161;102m█[0m[38;2;88;160;97m█[0m[38;2;117;163;103m█[0m[38;2;86;41;10m█[0m[38;2;250;202;95m█[0m[38;2;232;168;72m█[0m[38;2;236;176;83m█[0m[38;2;237;178;83m█[0m[38;2;239;177;81m█[0m[38;2;240;177;81m█[0m[38;2;238;177;83m█[0m[38;2;240;179;85m█[0m[38;2;239;176;83m█[0m[38;2;239;177;82m█[0m[38;2;245;182;93m█[0m[38;2;238;177;82m█[0m[38;2;238;177;83m█[0m[38;2;238;178;87m█[0m[38;2;238;176;79m█[0m[38;2;237;175;82m█[0m[38;2;239;176;81m█[0m[38;2;242;179;87m█[0m[38;2;135;88;35m█[0m[38;2;80;39;10m█[0m[38;2;246;220;197m█[0m[38;2;253;238;207m█[0m[38;2;255;239;207m█[0m[38;2;255;241;209m█[0m[38;2;252;239;207m█[0m[38;2;255;239;209m█[0m[38;2;156;121;88m█[0m[38;2;92;51;21m█[0m[38;2;183;159;119m█[0m[38;2;27;0;1m█[0m[38;2;142;112;79m█[0m[38;2;255;238;219m█[0m[38;2;254;241;209m█[0m[38;2;253;236;208m█[0m[38;2;255;239;210m█[0m[38;2;255;239;209m█[0m[38;2;253;237;206m█[0m[38;2;252;236;205m█[0m[38;2;255;238;209m█[0m[38;2;253;237;204m█[0m[38;2;253;236;208m█[0m[38;2;253;236;205m█[0m[38;2;254;237;209m█[0m[38;2;255;238;210m█[0m[38;2;253;238;207m█[0m[38;2;251;235;206m█[0m[38;2;75;37;13m█[0m[38;2;68;37;10m█[0m[38;2;255;239;200m█[0m[38;2;253;238;208m█[0m[38;2;254;239;208m█[0m[38;2;254;237;202m█[0m[38;2;47;19;5m█[0m[38;2;67;34;8m█[0m[38;2;70;35;6m█[0m[38;2;79;41;15m█[0m[38;2;72;37;9m█[0m[38;2;25;6;0m█[0m[38;2;242;179;88m█[0m[38;2;240;179;87m█[0m[38;2;240;181;89m█[0m[38;2;186;135;72m█[0m[38;2;76;39;9m█[0m[38;2;236;179;95m█[0m[38;2;241;181;90m█[0m[38;2;241;180;88m█[0m[38;2;236;180;84m█[0m[38;2;238;180;83m█[0m[38;2;239;178;86m█[0m[38;2;237;175;83m█[0m[38;2;236;174;81m█[0m[38;2;236;173;81m█[0m[38;2;240;179;86m█[0m[38;2;255;238;204m█[0m[38;2;231;181;93m█[0m[38;2;234;173;77m█[0m[38;2;233;173;79m█[0m[38;2;217;151;57m█[0m[38;2;79;47;15m█[0m[38;2;72;35;7m█[0m[38;2;75;153;109m█[0m[38;2;67;154;104m█[0m[38;2;63;151;106m█[0m[38;2;66;154;107m█[0m[38;2;66;150;96m█[0m[38;2;62;149;99m█[0m[38;2;61;146;100m█[0m");
$display("[38;2;137;182;60m█[0m[38;2;129;179;68m█[0m[38;2;153;192;55m█[0m[38;2;160;194;54m█[0m[38;2;160;194;47m█[0m[38;2;144;184;61m█[0m[38;2;160;192;52m█[0m[38;2;112;170;73m█[0m[38;2;129;181;69m█[0m[38;2;111;169;73m█[0m[38;2;155;189;56m█[0m[38;2;86;44;12m█[0m[38;2;65;17;2m█[0m[38;2;236;177;82m█[0m[38;2;238;179;84m█[0m[38;2;234;173;80m█[0m[38;2;240;175;83m█[0m[38;2;239;176;85m█[0m[38;2;236;177;81m█[0m[38;2;240;177;83m█[0m[38;2;237;179;85m█[0m[38;2;241;181;88m█[0m[38;2;239;179;84m█[0m[38;2;237;175;79m█[0m[38;2;239;179;86m█[0m[38;2;238;176;81m█[0m[38;2;238;178;88m█[0m[38;2;237;173;81m█[0m[38;2;242;178;84m█[0m[38;2;232;172;77m█[0m[38;2;236;174;81m█[0m[38;2;236;174;82m█[0m[38;2;60;20;0m█[0m[38;2;82;41;13m█[0m[38;2;254;238;208m█[0m[38;2;125;102;59m█[0m[38;2;79;40;11m█[0m[38;2;84;40;11m█[0m[38;2;84;44;14m█[0m[38;2;84;46;10m█[0m[38;2;47;8;0m█[0m[38;2;247;231;207m█[0m[38;2;253;254;246m█[0m[38;2;236;214;185m█[0m[38;2;92;52;23m█[0m[38;2;79;42;14m█[0m[38;2;80;42;13m█[0m[38;2;252;255;255m█[0m[38;2;253;237;205m█[0m[38;2;253;238;208m█[0m[38;2;252;238;204m█[0m[38;2;253;236;206m█[0m[38;2;253;237;205m█[0m[38;2;255;238;209m█[0m[38;2;253;237;205m█[0m[38;2;255;242;210m█[0m[38;2;254;239;206m█[0m[38;2;253;237;205m█[0m[38;2;255;237;208m█[0m[38;2;252;235;202m█[0m[38;2;83;42;15m█[0m[38;2;70;35;8m█[0m[38;2;75;38;13m█[0m[38;2;76;39;15m█[0m[38;2;72;38;14m█[0m[38;2;76;43;16m█[0m[38;2;254;238;207m█[0m[38;2;255;237;204m█[0m[38;2;253;239;209m█[0m[38;2;252;239;204m█[0m[38;2;254;237;211m█[0m[38;2;247;235;216m█[0m[38;2;236;174;82m█[0m[38;2;239;180;86m█[0m[38;2;233;171;76m█[0m[38;2;73;38;9m█[0m[38;2;77;43;12m█[0m[38;2;68;38;17m█[0m[38;2;246;184;87m█[0m[38;2;239;179;86m█[0m[38;2;237;177;81m█[0m[38;2;241;185;93m█[0m[38;2;233;175;81m█[0m[38;2;237;178;85m█[0m[38;2;238;179;82m█[0m[38;2;232;170;79m█[0m[38;2;234;172;78m█[0m[38;2;231;171;76m█[0m[38;2;210;145;50m█[0m[38;2;218;149;42m█[0m[38;2;79;37;9m█[0m[38;2;75;42;9m█[0m[38;2;122;173;72m█[0m[38;2;95;164;84m█[0m[38;2;99;165;82m█[0m[38;2;85;159;88m█[0m[38;2;111;171;69m█[0m[38;2;79;156;94m█[0m[38;2;81;158;87m█[0m[38;2;68;148;95m█[0m");
$display("[38;2;175;199;46m█[0m[38;2;159;189;41m█[0m[38;2;167;193;39m█[0m[38;2;173;200;50m█[0m[38;2;170;197;43m█[0m[38;2;180;202;38m█[0m[38;2;188;207;41m█[0m[38;2;180;203;40m█[0m[38;2;180;204;46m█[0m[38;2;180;205;42m█[0m[38;2;76;72;0m█[0m[38;2;88;46;14m█[0m[38;2;234;179;92m█[0m[38;2;238;179;85m█[0m[38;2;238;179;84m█[0m[38;2;237;176;81m█[0m[38;2;239;178;85m█[0m[38;2;240;177;86m█[0m[38;2;236;176;83m█[0m[38;2;239;178;86m█[0m[38;2;233;175;80m█[0m[38;2;239;176;82m█[0m[38;2;240;178;85m█[0m[38;2;236;179;84m█[0m[38;2;240;177;85m█[0m[38;2;236;174;81m█[0m[38;2;234;173;80m█[0m[38;2;237;173;79m█[0m[38;2;238;177;83m█[0m[38;2;236;177;78m█[0m[38;2;237;178;83m█[0m[38;2;236;174;81m█[0m[38;2;50;9;0m█[0m[38;2;87;47;13m█[0m[38;2;87;45;16m█[0m[38;2;255;252;240m█[0m[38;2;254;240;210m█[0m[38;2;254;240;208m█[0m[38;2;255;237;209m█[0m[38;2;254;239;208m█[0m[38;2;254;237;206m█[0m[38;2;253;237;205m█[0m[38;2;254;239;210m█[0m[38;2;254;238;208m█[0m[38;2;254;236;207m█[0m[38;2;255;240;211m█[0m[38;2;253;254;244m█[0m[38;2;85;47;21m█[0m[38;2;31;8;2m█[0m[38;2;254;239;208m█[0m[38;2;253;237;204m█[0m[38;2;255;239;209m█[0m[38;2;253;239;205m█[0m[38;2;254;235;204m█[0m[38;2;253;236;204m█[0m[38;2;254;235;204m█[0m[38;2;254;237;208m█[0m[38;2;254;238;205m█[0m[38;2;253;236;206m█[0m[38;2;252;235;205m█[0m[38;2;76;38;15m█[0m[38;2;84;54;28m█[0m[38;2;245;144;102m█[0m[38;2;244;147;108m█[0m[38;2;244;150;106m█[0m[38;2;78;42;15m█[0m[38;2;74;39;12m█[0m[38;2;255;239;207m█[0m[38;2;253;238;205m█[0m[38;2;255;239;210m█[0m[38;2;254;236;205m█[0m[38;2;253;236;206m█[0m[38;2;254;237;206m█[0m[38;2;234;176;76m█[0m[38;2;236;178;85m█[0m[38;2;239;177;84m█[0m[38;2;237;172;81m█[0m[38;2;226;170;73m█[0m[38;2;194;139;65m█[0m[38;2;236;176;82m█[0m[38;2;236;180;84m█[0m[38;2;237;175;82m█[0m[38;2;236;175;80m█[0m[38;2;234;173;80m█[0m[38;2;232;173;78m█[0m[38;2;81;32;0m█[0m[38;2;74;39;4m█[0m[38;2;219;147;38m█[0m[38;2;73;38;5m█[0m[38;2;78;41;8m█[0m[38;2;146;187;39m█[0m[38;2;136;179;47m█[0m[38;2;117;171;55m█[0m[38;2;148;185;44m█[0m[38;2;128;179;63m█[0m[38;2;149;187;41m█[0m[38;2;99;165;62m█[0m[38;2;109;167;56m█[0m[38;2;112;167;54m█[0m[38;2;79;150;77m█[0m");
$display("[38;2;174;195;38m█[0m[38;2;181;200;39m█[0m[38;2;192;204;40m█[0m[38;2;177;198;39m█[0m[38;2;182;201;40m█[0m[38;2;181;203;38m█[0m[38;2;170;194;32m█[0m[38;2;176;201;39m█[0m[38;2;175;199;38m█[0m[38;2;163;196;24m█[0m[38;2;87;40;6m█[0m[38;2;86;44;8m█[0m[38;2;236;175;74m█[0m[38;2;235;175;80m█[0m[38;2;241;181;86m█[0m[38;2;240;179;83m█[0m[38;2;237;177;83m█[0m[38;2;238;176;81m█[0m[38;2;240;179;82m█[0m[38;2;236;177;79m█[0m[38;2;238;179;86m█[0m[38;2;238;175;82m█[0m[38;2;237;173;80m█[0m[38;2;236;177;84m█[0m[38;2;237;179;83m█[0m[38;2;237;175;81m█[0m[38;2;238;177;86m█[0m[38;2;237;179;85m█[0m[38;2;240;180;87m█[0m[38;2;234;173;78m█[0m[38;2;232;171;77m█[0m[38;2;204;150;81m█[0m[38;2;85;44;10m█[0m[38;2;255;242;208m█[0m[38;2;254;238;206m█[0m[38;2;255;238;206m█[0m[38;2;253;238;205m█[0m[38;2;252;234;207m█[0m[38;2;255;238;207m█[0m[38;2;252;237;208m█[0m[38;2;254;238;209m█[0m[38;2;255;240;210m█[0m[38;2;254;239;206m█[0m[38;2;254;238;206m█[0m[38;2;254;237;209m█[0m[38;2;254;240;209m█[0m[38;2;254;239;207m█[0m[38;2;85;46;19m█[0m[38;2;78;42;11m█[0m[38;2;251;238;208m█[0m[38;2;253;237;206m█[0m[38;2;254;237;207m█[0m[38;2;253;237;205m█[0m[38;2;254;236;205m█[0m[38;2;251;234;203m█[0m[38;2;252;237;206m█[0m[38;2;252;235;203m█[0m[38;2;253;237;206m█[0m[38;2;254;237;204m█[0m[38;2;253;238;208m█[0m[38;2;248;255;254m█[0m[38;2;78;41;14m█[0m[38;2;255;118;65m█[0m[38;2;239;133;92m█[0m[38;2;237;132;91m█[0m[38;2;231;137;95m█[0m[38;2;78;44;14m█[0m[38;2;76;43;17m█[0m[38;2;249;239;220m█[0m[38;2;253;238;209m█[0m[38;2;250;234;203m█[0m[38;2;252;234;203m█[0m[38;2;255;237;206m█[0m[38;2;254;237;206m█[0m[38;2;251;239;209m█[0m[38;2;244;181;84m█[0m[38;2;237;178;85m█[0m[38;2;238;178;83m█[0m[38;2;238;176;81m█[0m[38;2;237;176;82m█[0m[38;2;234;176;80m█[0m[38;2;238;176;84m█[0m[38;2;237;176;83m█[0m[38;2;235;175;81m█[0m[38;2;204;142;45m█[0m[38;2;84;49;18m█[0m[38;2;81;44;11m█[0m[38;2;83;36;17m█[0m[38;2;154;195;31m█[0m[38;2;160;190;35m█[0m[38;2;154;187;37m█[0m[38;2;143;179;38m█[0m[38;2;145;183;44m█[0m[38;2;144;180;35m█[0m[38;2;153;186;41m█[0m[38;2;150;185;36m█[0m[38;2;140;178;38m█[0m[38;2;138;179;39m█[0m[38;2;139;178;36m█[0m[38;2;141;179;37m█[0m");
$display("[38;2;178;197;37m█[0m[38;2;206;209;46m█[0m[38;2;179;196;37m█[0m[38;2;217;214;50m█[0m[38;2;172;197;32m█[0m[38;2;167;193;32m█[0m[38;2;165;189;34m█[0m[38;2;75;29;7m█[0m[38;2;88;45;8m█[0m[38;2;101;57;18m█[0m[38;2;78;40;6m█[0m[38;2;87;43;6m█[0m[38;2;238;173;92m█[0m[38;2;236;178;84m█[0m[38;2;237;177;86m█[0m[38;2;236;176;83m█[0m[38;2;235;178;81m█[0m[38;2;236;174;81m█[0m[38;2;240;179;85m█[0m[38;2;236;175;84m█[0m[38;2;236;177;83m█[0m[38;2;240;178;86m█[0m[38;2;236;176;82m█[0m[38;2;238;178;82m█[0m[38;2;238;178;84m█[0m[38;2;236;173;79m█[0m[38;2;236;172;82m█[0m[38;2;235;175;80m█[0m[38;2;236;173;82m█[0m[38;2;239;178;84m█[0m[38;2;238;180;93m█[0m[38;2;84;43;12m█[0m[38;2;125;97;69m█[0m[38;2;255;238;209m█[0m[38;2;255;240;210m█[0m[38;2;254;236;206m█[0m[38;2;252;237;203m█[0m[38;2;254;238;207m█[0m[38;2;253;239;207m█[0m[38;2;253;239;210m█[0m[38;2;253;237;205m█[0m[38;2;253;239;207m█[0m[38;2;254;240;209m█[0m[38;2;246;231;200m█[0m[38;2;245;228;201m█[0m[38;2;254;238;206m█[0m[38;2;254;240;207m█[0m[38;2;84;44;15m█[0m[38;2;97;43;18m█[0m[38;2;254;237;209m█[0m[38;2;254;237;206m█[0m[38;2;252;236;206m█[0m[38;2;255;241;209m█[0m[38;2;255;236;203m█[0m[38;2;254;237;207m█[0m[38;2;255;237;206m█[0m[38;2;253;237;205m█[0m[38;2;252;235;200m█[0m[38;2;253;237;204m█[0m[38;2;253;235;205m█[0m[38;2;254;236;200m█[0m[38;2;255;241;206m█[0m[38;2;81;185;200m█[0m[38;2;78;92;80m█[0m[38;2;70;38;13m█[0m[38;2;81;44;16m█[0m[38;2;255;255;240m█[0m[38;2;246;241;202m█[0m[38;2;81;47;18m█[0m[38;2;68;35;8m█[0m[38;2;76;38;14m█[0m[38;2;255;242;210m█[0m[38;2;253;236;204m█[0m[38;2;254;238;206m█[0m[38;2;254;237;208m█[0m[38;2;244;129;90m█[0m[38;2;243;138;100m█[0m[38;2;242;130;90m█[0m[38;2;246;125;84m█[0m[38;2;242;118;82m█[0m[38;2;232;174;78m█[0m[38;2;237;176;81m█[0m[38;2;235;172;78m█[0m[38;2;208;145;52m█[0m[38;2;210;148;58m█[0m[38;2;68;35;11m█[0m[38;2;48;19;1m█[0m[38;2;152;179;31m█[0m[38;2;152;180;38m█[0m[38;2;178;191;41m█[0m[38;2;189;199;47m█[0m[38;2;155;186;39m█[0m[38;2;148;178;34m█[0m[38;2;156;186;39m█[0m[38;2;147;181;41m█[0m[38;2;147;183;35m█[0m[38;2;150;181;38m█[0m[38;2;127;169;30m█[0m[38;2;136;179;37m█[0m[38;2;149;185;47m█[0m");
$display("[38;2;201;205;45m█[0m[38;2;184;195;37m█[0m[38;2;191;200;42m█[0m[38;2;185;198;37m█[0m[38;2;166;194;39m█[0m[38;2;65;24;1m█[0m[38;2;84;43;6m█[0m[38;2;87;34;2m█[0m[38;2;252;237;207m█[0m[38;2;254;237;207m█[0m[38;2;254;238;207m█[0m[38;2;254;239;209m█[0m[38;2;253;238;206m█[0m[38;2;232;175;86m█[0m[38;2;236;178;84m█[0m[38;2;235;174;80m█[0m[38;2;237;177;83m█[0m[38;2;241;177;85m█[0m[38;2;240;179;86m█[0m[38;2;237;177;81m█[0m[38;2;239;179;85m█[0m[38;2;238;180;86m█[0m[38;2;242;178;86m█[0m[38;2;237;173;79m█[0m[38;2;237;176;83m█[0m[38;2;243;184;92m█[0m[38;2;238;178;87m█[0m[38;2;238;179;84m█[0m[38;2;235;176;82m█[0m[38;2;236;174;79m█[0m[38;2;255;213;109m█[0m[38;2;80;37;7m█[0m[38;2;250;237;206m█[0m[38;2;251;236;204m█[0m[38;2;255;241;209m█[0m[38;2;255;238;206m█[0m[38;2;253;238;206m█[0m[38;2;254;240;209m█[0m[38;2;254;236;207m█[0m[38;2;254;238;206m█[0m[38;2;255;238;208m█[0m[38;2;251;235;202m█[0m[38;2;252;235;202m█[0m[38;2;255;255;244m█[0m[38;2;243;233;213m█[0m[38;2;97;53;25m█[0m[38;2;84;42;14m█[0m[38;2;83;41;12m█[0m[38;2;252;236;205m█[0m[38;2;255;237;203m█[0m[38;2;253;236;204m█[0m[38;2;255;236;205m█[0m[38;2;253;238;204m█[0m[38;2;253;233;201m█[0m[38;2;254;236;202m██[0m[38;2;254;234;202m█[0m[38;2;253;235;205m█[0m[38;2;255;237;205m█[0m[38;2;252;236;202m█[0m[38;2;253;236;205m█[0m[38;2;253;236;204m█[0m[38;2;85;187;197m█[0m[38;2;255;231;197m█[0m[38;2;253;236;205m█[0m[38;2;254;238;207m█[0m[38;2;253;237;207m█[0m[38;2;253;239;207m█[0m[38;2;253;236;203m█[0m[38;2;255;235;205m█[0m[38;2;254;236;207m█[0m[38;2;254;236;204m█[0m[38;2;252;239;207m█[0m[38;2;254;237;205m█[0m[38;2;253;236;206m█[0m[38;2;246;140;102m█[0m[38;2;242;136;95m█[0m[38;2;247;146;105m█[0m[38;2;244;137;100m█[0m[38;2;255;243;214m█[0m[38;2;248;129;93m█[0m[38;2;246;180;93m█[0m[38;2;210;147;57m█[0m[38;2;206;142;51m█[0m[38;2;49;10;2m█[0m[38;2;78;42;15m█[0m[38;2;151;182;48m█[0m[38;2;137;173;33m█[0m[38;2;186;192;36m█[0m[38;2;196;201;46m█[0m[38;2;148;182;38m█[0m[38;2;180;198;43m█[0m[38;2;136;172;28m█[0m[38;2;161;184;35m█[0m[38;2;166;188;41m█[0m[38;2;148;179;35m█[0m[38;2;143;178;35m█[0m[38;2;146;181;36m█[0m[38;2;137;177;37m█[0m[38;2;149;181;37m█[0m");
$display("[38;2;167;191;39m█[0m[38;2;159;186;40m█[0m[38;2;160;189;37m█[0m[38;2;161;190;37m█[0m[38;2;82;45;12m█[0m[38;2;89;49;9m█[0m[38;2;250;235;208m█[0m[38;2;254;236;205m█[0m[38;2;253;237;205m█[0m[38;2;255;239;208m█[0m[38;2;255;240;208m█[0m[38;2;253;237;205m█[0m[38;2;254;236;206m█[0m[38;2;254;240;208m█[0m[38;2;253;237;206m█[0m[38;2;255;238;203m█[0m[38;2;248;233;212m█[0m[38;2;255;231;188m█[0m[38;2;220;165;72m█[0m[38;2;243;177;70m█[0m[38;2;243;180;77m█[0m[38;2;242;179;76m█[0m[38;2;225;163;74m█[0m[38;2;228;191;132m█[0m[38;2;252;250;219m█[0m[38;2;252;238;214m█[0m[38;2;254;238;203m█[0m[38;2;252;238;214m█[0m[38;2;255;237;206m█[0m[38;2;253;235;204m█[0m[38;2;127;100;71m█[0m[38;2;84;45;14m█[0m[38;2;254;242;207m█[0m[38;2;254;238;209m█[0m[38;2;253;236;204m█[0m[38;2;253;236;205m█[0m[38;2;254;238;206m█[0m[38;2;252;239;206m█[0m[38;2;254;236;203m█[0m[38;2;254;236;205m█[0m[38;2;254;237;206m█[0m[38;2;253;237;205m█[0m[38;2;252;239;206m█[0m[38;2;251;233;201m█[0m[38;2;254;236;204m█[0m[38;2;253;237;205m█[0m[38;2;253;234;202m█[0m[38;2;90;50;19m█[0m[38;2;83;44;16m█[0m[38;2;251;233;200m█[0m[38;2;253;236;202m█[0m[38;2;253;232;200m█[0m[38;2;253;238;206m█[0m[38;2;253;235;204m█[0m[38;2;251;233;201m█[0m[38;2;255;235;206m█[0m[38;2;253;237;207m█[0m[38;2;254;235;202m█[0m[38;2;253;236;205m█[0m[38;2;252;236;204m█[0m[38;2;252;236;205m█[0m[38;2;255;235;202m█[0m[38;2;92;179;186m█[0m[38;2;254;238;208m█[0m[38;2;253;236;206m█[0m[38;2;252;237;209m█[0m[38;2;254;238;208m█[0m[38;2;254;237;206m█[0m[38;2;251;233;203m█[0m[38;2;252;235;205m█[0m[38;2;252;235;204m█[0m[38;2;255;238;208m█[0m[38;2;255;238;209m█[0m[38;2;254;236;205m█[0m[38;2;253;238;206m█[0m[38;2;204;95;57m█[0m[38;2;243;134;95m█[0m[38;2;237;132;92m█[0m[38;2;240;138;101m█[0m[38;2;245;127;89m█[0m[38;2;244;123;84m█[0m[38;2;241;127;88m█[0m[38;2;233;204;162m█[0m[38;2;208;140;51m█[0m[38;2;72;41;11m█[0m[38;2;35;10;0m█[0m[38;2;138;173;38m█[0m[38;2;139;178;35m█[0m[38;2;151;176;30m█[0m[38;2;142;178;32m█[0m[38;2;157;184;38m█[0m[38;2;137;176;38m█[0m[38;2;158;186;42m█[0m[38;2;138;179;40m█[0m[38;2;142;177;40m█[0m[38;2;142;178;37m█[0m[38;2;136;172;34m█[0m[38;2;146;178;37m█[0m[38;2;147;179;38m█[0m[38;2;146;181;40m█[0m");
$display("[38;2;142;175;36m█[0m[38;2;148;180;39m█[0m[38;2;149;185;40m█[0m[38;2;94;100;10m█[0m[38;2;87;44;7m█[0m[38;2;254;235;202m█[0m[38;2;254;235;204m█[0m[38;2;253;236;207m█[0m[38;2;254;235;203m█[0m[38;2;253;237;208m█[0m[38;2;251;234;205m█[0m[38;2;254;237;207m█[0m[38;2;255;238;208m█[0m[38;2;254;237;207m█[0m[38;2;253;236;205m█[0m[38;2;254;238;205m█[0m[38;2;254;238;206m█[0m[38;2;253;237;207m█[0m[38;2;252;239;206m█[0m[38;2;253;236;203m█[0m[38;2;254;236;202m█[0m[38;2;253;233;203m█[0m[38;2;253;237;204m█[0m[38;2;253;235;205m█[0m[38;2;252;235;203m█[0m[38;2;253;237;206m█[0m[38;2;255;237;208m█[0m[38;2;252;236;208m█[0m[38;2;254;237;205m█[0m[38;2;252;236;204m█[0m[38;2;251;255;248m█[0m[38;2;71;36;12m█[0m[38;2;253;237;207m█[0m[38;2;255;239;210m█[0m[38;2;253;238;207m█[0m[38;2;253;236;209m█[0m[38;2;254;240;207m█[0m[38;2;254;237;206m█[0m[38;2;254;237;204m█[0m[38;2;255;238;208m█[0m[38;2;253;237;208m█[0m[38;2;253;238;210m█[0m[38;2;253;239;207m█[0m[38;2;254;239;209m█[0m[38;2;255;238;206m█[0m[38;2;253;236;202m█[0m[38;2;255;239;206m█[0m[38;2;80;41;12m█[0m[38;2;80;43;16m█[0m[38;2;229;201;161m█[0m[38;2;229;202;160m█[0m[38;2;254;235;204m█[0m[38;2;252;236;201m█[0m[38;2;254;233;199m█[0m[38;2;254;236;200m█[0m[38;2;251;234;199m█[0m[38;2;252;234;204m█[0m[38;2;253;237;203m█[0m[38;2;252;236;200m█[0m[38;2;253;236;203m█[0m[38;2;251;236;206m█[0m[38;2;238;250;228m█[0m[38;2;60;188;207m█[0m[38;2;253;237;207m█[0m[38;2;253;238;208m█[0m[38;2;255;236;206m█[0m[38;2;253;236;203m█[0m[38;2;253;235;201m█[0m[38;2;254;237;205m█[0m[38;2;254;236;205m█[0m[38;2;253;236;203m█[0m[38;2;254;239;205m█[0m[38;2;252;238;206m█[0m[38;2;253;240;206m█[0m[38;2;253;237;206m█[0m[38;2;252;240;206m█[0m[38;2;248;241;208m█[0m[38;2;242;113;74m█[0m[38;2;241;132;96m█[0m[38;2;239;120;83m█[0m[38;2;240;129;92m█[0m[38;2;244;214;177m█[0m[38;2;229;205;163m█[0m[38;2;64;32;5m█[0m[38;2;54;40;5m█[0m[38;2;82;143;41m█[0m[38;2;62;129;26m█[0m[38;2;107;160;35m█[0m[38;2;112;160;36m█[0m[38;2;104;158;37m█[0m[38;2;115;168;42m█[0m[38;2;113;165;41m█[0m[38;2;115;167;38m█[0m[38;2;116;166;38m█[0m[38;2;125;169;39m█[0m[38;2;116;163;37m█[0m[38;2;122;165;37m█[0m[38;2;118;165;38m█[0m[38;2;129;169;35m█[0m[38;2;121;165;37m█[0m");
$display("[38;2;152;183;39m█[0m[38;2;145;178;37m█[0m[38;2;134;173;34m█[0m[38;2;46;34;1m█[0m[38;2;81;43;10m█[0m[38;2;252;240;205m█[0m[38;2;254;237;206m█[0m[38;2;253;244;205m█[0m[38;2;30;6;0m█[0m[38;2;255;238;205m█[0m[38;2;255;237;207m█[0m[38;2;252;237;206m█[0m[38;2;254;236;202m█[0m[38;2;252;236;207m█[0m[38;2;255;238;207m█[0m[38;2;254;237;206m█[0m[38;2;252;236;206m█[0m[38;2;255;238;209m█[0m[38;2;253;237;206m█[0m[38;2;254;237;207m█[0m[38;2;253;236;206m█[0m[38;2;253;236;203m█[0m[38;2;253;234;202m█[0m[38;2;254;239;206m█[0m[38;2;252;235;204m█[0m[38;2;255;239;209m█[0m[38;2;255;235;206m█[0m[38;2;254;238;207m█[0m[38;2;255;237;205m█[0m[38;2;253;234;204m█[0m[38;2;254;235;201m█[0m[38;2;72;38;13m█[0m[38;2;72;32;8m█[0m[38;2;254;238;209m██[0m[38;2;255;235;205m█[0m[38;2;255;236;206m█[0m[38;2;253;236;206m█[0m[38;2;254;237;204m█[0m[38;2;254;236;202m█[0m[38;2;253;237;206m█[0m[38;2;254;238;204m█[0m[38;2;253;237;203m█[0m[38;2;252;237;205m█[0m[38;2;255;237;207m█[0m[38;2;252;236;204m█[0m[38;2;239;210;173m█[0m[38;2;66;34;9m█[0m[38;2;34;7;0m█[0m[38;2;228;201;158m█[0m[38;2;227;197;152m█[0m[38;2;227;198;155m█[0m[38;2;229;199;158m█[0m[38;2;228;198;156m█[0m[38;2;255;241;205m█[0m[38;2;254;238;202m█[0m[38;2;253;232;200m█[0m[38;2;253;235;204m█[0m[38;2;254;235;201m█[0m[38;2;249;233;197m█[0m[38;2;253;234;204m█[0m[38;2;251;237;206m█[0m[38;2;90;194;200m█[0m[38;2;250;231;203m█[0m[38;2;254;235;198m█[0m[38;2;255;235;204m█[0m[38;2;252;235;204m█[0m[38;2;252;232;200m█[0m[38;2;252;235;203m█[0m[38;2;253;237;205m█[0m[38;2;253;235;203m█[0m[38;2;254;238;209m█[0m[38;2;254;236;204m█[0m[38;2;253;237;202m█[0m[38;2;254;234;205m█[0m[38;2;253;236;203m█[0m[38;2;255;238;206m█[0m[38;2;232;209;167m█[0m[38;2;231;204;168m█[0m[38;2;230;203;163m█[0m[38;2;229;202;165m█[0m[38;2;228;202;158m█[0m[38;2;226;201;156m█[0m[38;2;57;30;7m█[0m[38;2;37;22;0m█[0m[38;2;49;119;49m█[0m[38;2;37;109;39m█[0m[38;2;41;113;39m█[0m[38;2;85;149;46m█[0m[38;2;37;113;45m█[0m[38;2;54;124;36m█[0m[38;2;85;146;42m█[0m[38;2;95;156;38m█[0m[38;2;95;154;41m█[0m[38;2;95;151;35m█[0m[38;2;80;146;37m█[0m[38;2;95;153;38m█[0m[38;2;102;156;41m█[0m[38;2;96;152;36m█[0m[38;2;105;158;39m█[0m");
$display("[38;2;118;167;39m█[0m[38;2;124;169;33m█[0m[38;2;120;167;41m█[0m[38;2;118;168;36m█[0m[38;2;67;42;9m█[0m[38;2;74;40;11m█[0m[38;2;19;1;2m█[0m[38;2;72;39;10m█[0m[38;2;252;239;200m█[0m[38;2;252;229;186m█[0m[38;2;253;240;213m█[0m[38;2;253;241;211m█[0m[38;2;241;211;173m█[0m[38;2;228;205;164m█[0m[38;2;231;206;167m█[0m[38;2;234;210;169m█[0m[38;2;237;209;167m█[0m[38;2;229;200;162m█[0m[38;2;235;208;169m█[0m[38;2;229;204;167m█[0m[38;2;248;237;207m█[0m[38;2;255;235;201m█[0m[38;2;255;238;205m█[0m[38;2;250;238;202m█[0m[38;2;252;237;205m█[0m[38;2;253;235;204m█[0m[38;2;253;236;204m█[0m[38;2;253;236;203m█[0m[38;2;253;238;207m█[0m[38;2;254;239;205m█[0m[38;2;254;239;206m█[0m[38;2;16;0;0m█[0m[38;2;66;36;10m█[0m[38;2;250;237;196m█[0m[38;2;254;236;204m█[0m[38;2;253;236;202m█[0m[38;2;250;234;201m█[0m[38;2;252;236;205m█[0m[38;2;252;236;204m█[0m[38;2;253;236;204m█[0m[38;2;254;238;207m█[0m[38;2;255;237;204m█[0m[38;2;254;237;203m█[0m[38;2;253;236;203m█[0m[38;2;250;241;210m█[0m[38;2;230;201;162m█[0m[38;2;67;38;15m█[0m[38;2;65;37;9m█[0m[38;2;222;192;152m█[0m[38;2;226;197;154m█[0m[38;2;216;188;145m█[0m[38;2;224;194;151m█[0m[38;2;222;195;149m█[0m[38;2;226;199;157m█[0m[38;2;219;188;142m█[0m[38;2;223;197;152m█[0m[38;2;222;193;148m█[0m[38;2;221;188;146m█[0m[38;2;228;195;152m█[0m[38;2;218;188;144m█[0m[38;2;252;238;204m█[0m[38;2;241;237;214m█[0m[38;2;112;200;199m█[0m[38;2;110;204;204m█[0m[38;2;47;176;196m█[0m[38;2;245;237;212m█[0m[38;2;253;236;206m█[0m[38;2;250;234;205m█[0m[38;2;253;233;202m█[0m[38;2;254;234;199m█[0m[38;2;253;232;200m█[0m[38;2;252;237;202m█[0m[38;2;250;233;194m█[0m[38;2;230;206;166m█[0m[38;2;236;206;166m█[0m[38;2;231;207;166m█[0m[38;2;232;204;165m█[0m[38;2;224;197;157m█[0m[38;2;227;202;162m█[0m[38;2;231;205;162m█[0m[38;2;231;205;166m█[0m[38;2;73;35;15m█[0m[38;2;58;36;9m█[0m[38;2;50;24;3m█[0m[38;2;30;102;44m█[0m[38;2;23;94;39m█[0m[38;2;33;103;46m█[0m[38;2;27;98;40m█[0m[38;2;36;108;45m█[0m[38;2;45;119;46m█[0m[38;2;55;125;48m█[0m[38;2;41;113;43m█[0m[38;2;66;135;51m█[0m[38;2;54;125;45m█[0m[38;2;61;128;44m█[0m[38;2;75;143;43m█[0m[38;2;53;130;47m█[0m[38;2;75;142;36m█[0m[38;2;90;150;39m█[0m[38;2;95;156;44m█[0m");
$display("[38;2;114;163;41m█[0m[38;2;112;159;39m█[0m[38;2;77;139;38m█[0m[38;2;78;140;45m█[0m[38;2;75;139;50m█[0m[38;2;57;121;40m█[0m[38;2;66;70;23m█[0m[38;2;67;36;9m█[0m[38;2;70;38;11m█[0m[38;2;70;36;7m█[0m[38;2;71;38;12m█[0m[38;2;70;37;7m█[0m[38;2;73;38;16m█[0m[38;2;66;38;11m█[0m[38;2;65;37;12m█[0m[38;2;62;33;9m█[0m[38;2;67;30;7m█[0m[38;2;64;34;10m█[0m[38;2;69;40;15m█[0m[38;2;69;38;9m█[0m[38;2;70;39;10m█[0m[38;2;63;32;5m█[0m[38;2;63;35;13m█[0m[38;2;41;16;0m█[0m[38;2;252;239;200m█[0m[38;2;242;219;181m█[0m[38;2;225;198;154m█[0m[38;2;224;199;154m█[0m[38;2;229;201;158m█[0m[38;2;229;202;159m█[0m[38;2;226;198;156m█[0m[38;2;255;240;202m█[0m[38;2;50;23;2m█[0m[38;2;66;38;10m█[0m[38;2;71;39;11m█[0m[38;2;235;214;173m█[0m[38;2;231;205;167m█[0m[38;2;235;210;171m█[0m[38;2;236;210;172m█[0m[38;2;232;207;169m█[0m[38;2;228;202;162m█[0m[38;2;228;202;164m█[0m[38;2;229;203;166m█[0m[38;2;232;207;163m█[0m[38;2;255;243;204m█[0m[38;2;65;36;9m█[0m[38;2;69;38;15m█[0m[38;2;53;94;45m█[0m[38;2;61;31;8m█[0m[38;2;55;27;3m█[0m[38;2;59;34;12m█[0m[38;2;62;39;10m█[0m[38;2;42;20;4m█[0m[38;2;219;189;142m█[0m[38;2;218;187;143m█[0m[38;2;224;194;145m█[0m[38;2;227;196;157m█[0m[38;2;111;173;160m█[0m[38;2;62;190;202m█[0m[38;2;74;195;215m█[0m[38;2;78;191;196m█[0m[38;2;126;216;216m█[0m[38;2;118;207;204m█[0m[38;2;122;210;208m█[0m[38;2;120;210;209m█[0m[38;2;121;208;206m█[0m[38;2;119;206;201m█[0m[38;2;119;207;206m█[0m[38;2;87;189;199m█[0m[38;2;227;202;156m█[0m[38;2;232;203;161m█[0m[38;2;229;204;163m█[0m[38;2;228;200;158m█[0m[38;2;224;199;154m█[0m[38;2;229;202;159m█[0m[38;2;231;201;159m█[0m[38;2;228;200;157m█[0m[38;2;244;229;194m█[0m[38;2;66;40;15m█[0m[38;2;60;35;11m█[0m[38;2;56;34;13m█[0m[38;2;62;32;12m█[0m[38;2;35;100;48m█[0m[38;2;29;98;44m█[0m[38;2;26;97;43m█[0m[38;2;20;89;34m█[0m[38;2;34;104;38m█[0m[38;2;37;110;47m█[0m[38;2;36;108;42m█[0m[38;2;37;107;42m█[0m[38;2;37;106;46m█[0m[38;2;50;121;36m█[0m[38;2;40;110;46m█[0m[38;2;41;115;44m█[0m[38;2;50;120;43m█[0m[38;2;54;128;41m█[0m[38;2;44;116;43m█[0m[38;2;46;117;43m█[0m[38;2;50;120;41m█[0m[38;2;62;130;40m█[0m");
$display("[38;2;107;159;40m█[0m[38;2;112;161;41m█[0m[38;2;104;155;38m█[0m[38;2;108;160;41m█[0m[38;2;85;145;32m█[0m[38;2;99;151;42m█[0m[38;2;73;132;45m█[0m[38;2;69;132;36m█[0m[38;2;67;129;39m█[0m[38;2;109;154;40m█[0m[38;2;107;152;41m█[0m[38;2;51;112;37m█[0m[38;2;56;120;49m█[0m[38;2;85;143;40m█[0m[38;2;60;124;46m█[0m[38;2;59;125;44m█[0m[38;2;50;114;34m█[0m[38;2;77;135;42m█[0m[38;2;51;120;42m█[0m[38;2;43;102;40m█[0m[38;2;41;105;41m█[0m[38;2;53;114;42m█[0m[38;2;40;110;29m█[0m[38;2;46;111;46m█[0m[38;2;66;84;41m█[0m[38;2;48;35;4m█[0m[38;2;47;24;0m█[0m[38;2;53;27;0m█[0m[38;2;55;29;0m█[0m[38;2;52;29;2m█[0m[38;2;36;18;0m█[0m[38;2;48;48;13m█[0m[38;2;43;110;46m█[0m[38;2;41;102;42m█[0m[38;2;65;125;53m█[0m[38;2;67;37;11m█[0m[38;2;66;36;9m█[0m[38;2;70;40;11m█[0m[38;2;66;36;8m█[0m[38;2;66;38;12m█[0m[38;2;64;33;9m█[0m[38;2;66;38;10m█[0m[38;2;68;36;9m█[0m[38;2;55;33;1m█[0m[38;2;50;40;9m█[0m[38;2;40;105;38m█[0m[38;2;43;104;37m█[0m[38;2;40;106;37m█[0m[38;2;50;118;45m█[0m[38;2;34;97;39m█[0m[38;2;43;111;42m█[0m[38;2;38;105;41m█[0m[38;2;53;102;48m█[0m[38;2;71;33;10m█[0m[38;2;87;185;195m█[0m[38;2;125;207;209m█[0m[38;2;194;229;224m█[0m[38;2;193;229;220m█[0m[38;2;110;208;215m█[0m[38;2;125;209;210m█[0m[38;2;129;211;213m█[0m[38;2;127;212;211m█[0m[38;2;124;210;207m█[0m[38;2;120;208;204m█[0m[38;2;118;206;205m█[0m[38;2;113;205;205m█[0m[38;2;114;204;206m█[0m[38;2;113;202;203m█[0m[38;2;122;211;210m█[0m[38;2;126;211;210m█[0m[38;2;89;186;193m█[0m[38;2;117;171;167m█[0m[38;2;56;35;10m█[0m[38;2;57;35;8m█[0m[38;2;53;32;6m█[0m[38;2;59;31;8m█[0m[38;2;61;30;6m█[0m[38;2;57;81;42m█[0m[38;2;21;92;36m█[0m[38;2;37;104;41m█[0m[38;2;34;102;41m█[0m[38;2;36;105;42m█[0m[38;2;33;103;39m█[0m[38;2;42;115;53m█[0m[38;2;63;133;41m█[0m[38;2;75;143;47m█[0m[38;2;37;110;43m█[0m[38;2;67;137;40m█[0m[38;2;82;147;47m█[0m[38;2;59;128;43m█[0m[38;2;53;124;37m█[0m[38;2;73;142;47m█[0m[38;2;42;115;38m█[0m[38;2;65;132;42m█[0m[38;2;68;139;50m█[0m[38;2;71;139;44m█[0m[38;2;58;127;46m█[0m[38;2;76;143;44m█[0m[38;2;81;148;44m█[0m[38;2;71;139;42m█[0m");
$display("[38;2;115;164;38m█[0m[38;2;117;162;39m█[0m[38;2;123;166;37m█[0m[38;2;119;163;40m█[0m[38;2;112;156;34m█[0m[38;2;113;159;37m█[0m[38;2;111;158;42m█[0m[38;2;105;154;31m█[0m[38;2;110;158;37m█[0m[38;2;101;152;37m█[0m[38;2;126;165;37m█[0m[38;2;134;173;40m█[0m[38;2;110;158;37m█[0m[38;2;114;162;38m█[0m[38;2;111;162;39m█[0m[38;2;82;142;33m█[0m[38;2;93;151;43m█[0m[38;2;84;143;35m█[0m[38;2;99;154;41m█[0m[38;2;95;150;40m█[0m[38;2;51;119;35m█[0m[38;2;103;155;40m█[0m[38;2;89;146;47m█[0m[38;2;101;151;37m█[0m[38;2;96;151;39m█[0m[38;2;101;154;38m█[0m[38;2;70;132;36m█[0m[38;2;66;130;38m█[0m[38;2;74;139;48m█[0m[38;2;60;123;38m█[0m[38;2;61;124;41m█[0m[38;2;75;129;37m█[0m[38;2;69;132;45m█[0m[38;2;74;136;49m█[0m[38;2;64;132;45m█[0m[38;2;60;124;35m█[0m[38;2;61;126;46m█[0m[38;2;59;124;41m█[0m[38;2;55;118;39m█[0m[38;2;46;115;36m█[0m[38;2;51;112;36m█[0m[38;2;60;122;42m█[0m[38;2;52;120;43m█[0m[38;2;49;118;38m█[0m[38;2;41;106;34m█[0m[38;2;83;143;38m█[0m[38;2;57;123;42m█[0m[38;2;58;122;42m█[0m[38;2;55;125;36m█[0m[38;2;53;122;41m█[0m[38;2;61;127;44m█[0m[38;2;56;122;37m█[0m[38;2;57;121;41m█[0m[38;2;56;120;41m█[0m[38;2;82;184;190m█[0m[38;2;117;206;206m█[0m[38;2;123;206;206m█[0m[38;2;122;209;207m█[0m[38;2;121;207;207m█[0m[38;2;156;222;219m█[0m[38;2;170;231;228m█[0m[38;2;122;209;206m█[0m[38;2;119;208;205m█[0m[38;2;119;208;207m█[0m[38;2;163;230;228m█[0m[38;2;159;225;221m█[0m[38;2;112;206;206m█[0m[38;2;111;203;205m█[0m[38;2;115;209;208m█[0m[38;2;107;198;201m█[0m[38;2;119;210;210m█[0m[38;2;112;199;200m█[0m[38;2;75;179;199m█[0m[38;2;37;108;45m█[0m[38;2;41;109;42m█[0m[38;2;43;112;41m█[0m[38;2;61;126;41m█[0m[38;2;50;116;39m█[0m[38;2;61;131;50m█[0m[38;2;65;134;37m█[0m[38;2;75;142;44m█[0m[38;2;80;145;45m█[0m[38;2;48;118;52m█[0m[38;2;69;137;41m█[0m[38;2;73;140;44m█[0m[38;2;74;142;42m█[0m[38;2;82;147;40m█[0m[38;2;72;138;34m█[0m[38;2;81;148;43m█[0m[38;2;76;143;39m█[0m[38;2;73;141;43m█[0m[38;2;71;142;42m█[0m[38;2;76;144;42m█[0m[38;2;70;140;44m█[0m[38;2;68;141;46m█[0m[38;2;73;144;44m█[0m[38;2;68;138;37m█[0m[38;2;73;145;44m█[0m[38;2;65;140;39m█[0m[38;2;75;145;44m█[0m");
$display("[38;2;93;152;43m█[0m[38;2;105;157;37m█[0m[38;2;119;165;47m█[0m[38;2;112;158;35m█[0m[38;2;104;158;39m█[0m[38;2;102;151;32m█[0m[38;2;110;158;34m█[0m[38;2;109;159;39m█[0m[38;2;110;157;36m█[0m[38;2;156;178;38m█[0m[38;2;121;163;38m█[0m[38;2;114;163;35m█[0m[38;2;122;165;41m█[0m[38;2;124;165;38m█[0m[38;2;119;162;34m█[0m[38;2;120;162;37m█[0m[38;2;124;171;40m█[0m[38;2;117;162;39m█[0m[38;2;121;165;35m█[0m[38;2;120;164;32m█[0m[38;2;126;167;41m█[0m[38;2;103;154;34m█[0m[38;2;128;170;44m█[0m[38;2;124;167;38m█[0m[38;2;115;158;35m█[0m[38;2;118;165;39m█[0m[38;2;128;170;42m█[0m[38;2;108;160;35m█[0m[38;2;101;155;39m█[0m[38;2;106;159;38m█[0m[38;2;116;155;28m█[0m[38;2;119;165;40m█[0m[38;2;122;163;37m█[0m[38;2;122;167;40m█[0m[38;2;96;154;46m█[0m[38;2;127;170;44m█[0m[38;2;114;161;38m█[0m[38;2;85;145;44m█[0m[38;2;93;151;43m█[0m[38;2;104;157;43m█[0m[38;2;91;147;38m█[0m[38;2;84;146;50m█[0m[38;2;121;164;44m█[0m[38;2;77;136;37m█[0m[38;2;95;147;33m█[0m[38;2;116;165;41m█[0m[38;2;79;144;53m█[0m[38;2;109;159;41m█[0m[38;2;106;161;39m█[0m[38;2;79;137;37m█[0m[38;2;78;137;37m█[0m[38;2;87;148;48m█[0m[38;2;67;129;42m█[0m[38;2;74;138;46m█[0m[38;2;78;138;38m█[0m[38;2;72;135;45m█[0m[38;2;58;126;49m█[0m[38;2;44;115;39m█[0m[38;2;85;183;193m█[0m[38;2;109;200;203m█[0m[38;2;118;202;203m█[0m[38;2;118;206;208m█[0m[38;2;129;213;212m█[0m[38;2;130;210;208m█[0m[38;2;111;203;206m█[0m[38;2;105;196;200m█[0m[38;2;106;200;202m█[0m[38;2;106;198;199m█[0m[38;2;104;198;204m█[0m[38;2;85;192;214m█[0m[38;2;49;101;21m█[0m[38;2;39;111;49m█[0m[38;2;54;121;45m█[0m[38;2;45;119;47m█[0m[38;2;69;134;41m█[0m[38;2;56;128;49m█[0m[38;2;80;141;38m█[0m[38;2;72;141;39m█[0m[38;2;77;142;39m█[0m[38;2;77;142;41m█[0m[38;2;79;148;46m█[0m[38;2;88;149;41m█[0m[38;2;76;140;35m█[0m[38;2;81;146;42m█[0m[38;2;72;143;39m█[0m[38;2;69;138;43m█[0m[38;2;67;139;40m█[0m[38;2;74;141;39m█[0m[38;2;69;140;47m█[0m[38;2;74;144;44m█[0m[38;2;71;141;42m█[0m[38;2;58;131;39m█[0m[38;2;78;146;46m█[0m[38;2;72;142;44m█[0m[38;2;68;138;48m█[0m[38;2;72;142;44m█[0m[38;2;76;144;46m█[0m[38;2;68;143;51m█[0m[38;2;63;132;38m█[0m[38;2;65;135;43m█[0m");
$display("[38;2;90;151;44m█[0m[38;2;91;149;46m█[0m[38;2;87;149;42m█[0m[38;2;118;162;41m█[0m[38;2;142;172;40m█[0m[38;2;99;157;39m█[0m[38;2;95;151;39m█[0m[38;2;138;170;38m█[0m[38;2;111;161;42m█[0m[38;2;113;163;43m█[0m[38;2;161;183;45m█[0m[38;2;108;157;34m█[0m[38;2;113;161;40m█[0m[38;2;122;166;40m█[0m[38;2;109;159;38m█[0m[38;2;117;161;35m█[0m[38;2;104;155;38m█[0m[38;2;118;162;40m█[0m[38;2;122;167;41m█[0m[38;2;125;167;36m█[0m[38;2;121;165;40m█[0m[38;2;114;160;37m█[0m[38;2;126;163;31m█[0m[38;2;123;165;35m█[0m[38;2;139;173;39m█[0m[38;2;124;165;38m█[0m[38;2;119;160;35m█[0m[38;2;160;181;39m█[0m[38;2;155;182;42m█[0m[38;2;124;164;35m█[0m[38;2;123;166;38m█[0m[38;2;129;168;37m█[0m[38;2;127;168;39m█[0m[38;2;139;173;37m█[0m[38;2;131;168;32m█[0m[38;2;132;169;37m█[0m[38;2;130;171;40m█[0m[38;2;125;166;31m█[0m[38;2;129;169;41m█[0m[38;2;119;163;34m█[0m[38;2;118;159;30m█[0m[38;2;121;162;35m█[0m[38;2;122;164;32m█[0m[38;2;123;161;29m█[0m[38;2;126;164;32m█[0m[38;2;125;164;32m█[0m[38;2;132;172;38m█[0m[38;2;125;167;43m█[0m[38;2;122;166;37m█[0m[38;2;106;158;37m█[0m[38;2;117;161;33m█[0m[38;2;108;157;38m█[0m[38;2;114;160;38m█[0m[38;2;108;155;39m█[0m[38;2;102;153;38m█[0m[38;2;114;163;42m█[0m[38;2;100;155;40m█[0m[38;2;94;151;42m█[0m[38;2;92;150;39m█[0m[38;2;68;131;36m█[0m[38;2;68;140;38m█[0m[38;2;101;197;199m█[0m[38;2;62;174;199m█[0m[38;2;71;179;204m█[0m[38;2;70;179;195m█[0m[38;2;84;187;206m█[0m[38;2;43;126;89m█[0m[38;2;62;132;44m█[0m[38;2;54;121;37m█[0m[38;2;62;128;46m█[0m[38;2;52;122;36m█[0m[38;2;93;148;37m█[0m[38;2;91;150;43m█[0m[38;2;80;148;44m█[0m[38;2;77;142;37m█[0m[38;2;88;147;42m█[0m[38;2;103;158;45m█[0m[38;2;83;146;40m█[0m[38;2;80;145;39m█[0m[38;2;83;149;42m█[0m[38;2;82;147;40m█[0m[38;2;81;146;42m█[0m[38;2;80;145;40m█[0m[38;2;73;140;44m█[0m[38;2;71;140;42m█[0m[38;2;73;142;41m█[0m[38;2;80;147;43m█[0m[38;2;129;170;46m█[0m[38;2;71;142;40m█[0m[38;2;68;140;45m█[0m[38;2;75;144;44m█[0m[38;2;128;174;53m█[0m[38;2;130;175;57m█[0m[38;2;76;147;44m█[0m[38;2;70;145;48m█[0m[38;2;61;138;42m█[0m[38;2;55;130;47m█[0m[38;2;63;136;46m█[0m[38;2;55;131;40m█[0m[38;2;62;136;47m█[0m");
$display("[38;2;71;143;46m█[0m[38;2;73;137;41m█[0m[38;2;76;146;40m█[0m[38;2;78;144;41m█[0m[38;2;77;141;40m█[0m[38;2;123;166;41m█[0m[38;2;98;155;41m█[0m[38;2;79;143;35m█[0m[38;2;105;153;37m█[0m[38;2;96;154;43m█[0m[38;2;109;157;36m█[0m[38;2;128;169;41m█[0m[38;2;104;156;38m█[0m[38;2;97;149;34m█[0m[38;2;83;140;42m█[0m[38;2;73;142;45m█[0m[38;2;95;156;41m█[0m[38;2;108;159;38m█[0m[38;2;109;158;35m█[0m[38;2;105;154;36m█[0m[38;2;117;166;41m█[0m[38;2;117;163;39m█[0m[38;2;115;160;34m█[0m[38;2;116;164;35m█[0m[38;2;128;168;40m█[0m[38;2;149;177;40m█[0m[38;2;186;191;42m█[0m[38;2;169;194;50m█[0m[38;2;169;188;41m█[0m[38;2;160;183;41m█[0m[38;2;117;163;42m█[0m[38;2;125;168;35m█[0m[38;2;150;179;39m█[0m[38;2;147;182;46m█[0m[38;2;118;163;35m█[0m[38;2;117;159;35m█[0m[38;2;141;178;45m█[0m[38;2;131;169;33m█[0m[38;2;132;170;36m█[0m[38;2;125;165;34m█[0m[38;2;124;166;33m█[0m[38;2;125;168;36m█[0m[38;2;126;169;36m█[0m[38;2;125;171;38m█[0m[38;2;123;166;34m█[0m[38;2;123;165;33m█[0m[38;2;127;170;40m█[0m[38;2;120;164;38m█[0m[38;2;131;169;38m█[0m[38;2;132;173;42m█[0m[38;2;129;168;39m█[0m[38;2;130;167;37m█[0m[38;2;121;165;38m█[0m[38;2;113;158;34m█[0m[38;2;119;162;36m█[0m[38;2;120;162;38m█[0m[38;2;113;159;36m█[0m[38;2;109;161;39m█[0m[38;2;102;156;40m█[0m[38;2;96;149;36m█[0m[38;2;100;155;41m█[0m[38;2;98;152;41m█[0m[38;2;76;144;41m█[0m[38;2;82;144;40m█[0m[38;2;94;155;41m█[0m[38;2;104;155;36m█[0m[38;2;99;149;36m█[0m[38;2;90;151;45m█[0m[38;2;93;150;42m█[0m[38;2;93;150;39m█[0m[38;2;95;151;38m█[0m[38;2;96;152;37m█[0m[38;2;92;148;40m█[0m[38;2;87;149;41m█[0m[38;2;91;149;39m█[0m[38;2;91;149;40m█[0m[38;2;132;165;41m█[0m[38;2;122;167;44m█[0m[38;2;79;142;32m█[0m[38;2;88;152;44m█[0m[38;2;89;153;44m█[0m[38;2;75;140;41m█[0m[38;2;69;139;46m█[0m[38;2;67;135;46m█[0m[38;2;80;144;40m█[0m[38;2;91;152;45m█[0m[38;2;107;152;33m█[0m[38;2;69;140;39m█[0m[38;2;76;143;43m█[0m[38;2;125;164;44m█[0m[38;2;131;168;48m█[0m[38;2;77;144;42m█[0m[38;2;70;142;45m█[0m[38;2;73;146;47m█[0m[38;2;89;149;36m█[0m[38;2;69;143;47m█[0m[38;2;59;134;45m█[0m[38;2;67;141;51m█[0m[38;2;67;142;47m█[0m[38;2;54;132;46m█[0m");
$display("[38;2;49;121;51m█[0m[38;2;42;119;49m█[0m[38;2;56;127;49m█[0m[38;2;76;146;45m█[0m[38;2;72;141;42m█[0m[38;2;57;130;49m█[0m[38;2;58;125;46m█[0m[38;2;82;149;53m█[0m[38;2;72;141;41m█[0m[38;2;104;161;50m█[0m[38;2;85;147;44m█[0m[38;2;62;134;47m█[0m[38;2;91;151;48m█[0m[38;2;60;130;50m█[0m[38;2;56;130;44m█[0m[38;2;82;147;40m█[0m[38;2;93;150;40m█[0m[38;2;88;150;39m█[0m[38;2;69;136;42m█[0m[38;2;82;142;47m█[0m[38;2;102;157;45m█[0m[38;2;103;158;41m█[0m[38;2;112;162;39m█[0m[38;2;123;164;33m█[0m[38;2;124;166;38m█[0m[38;2;112;158;36m█[0m[38;2;119;161;38m█[0m[38;2;144;173;40m█[0m[38;2;150;182;51m█[0m[38;2;133;166;36m█[0m[38;2;142;173;35m█[0m[38;2;129;165;37m█[0m[38;2;146;175;37m█[0m[38;2;111;158;39m█[0m[38;2;135;164;31m█[0m[38;2;136;169;33m█[0m[38;2;112;162;39m█[0m[38;2;124;164;38m█[0m[38;2;115;158;34m█[0m[38;2;126;163;32m█[0m[38;2;123;164;37m█[0m[38;2;121;168;40m█[0m[38;2;116;163;40m█[0m[38;2;117;166;41m█[0m[38;2;131;170;39m█[0m[38;2;119;159;33m█[0m[38;2;123;164;38m█[0m[38;2;119;163;37m█[0m[38;2;122;167;42m█[0m[38;2;122;164;38m█[0m[38;2;120;161;35m█[0m[38;2;114;163;44m█[0m[38;2;119;164;39m█[0m[38;2;114;159;35m█[0m[38;2;108;160;44m█[0m[38;2;101;158;43m█[0m[38;2;108;159;39m█[0m[38;2;106;159;42m█[0m[38;2;93;151;37m█[0m[38;2;93;149;36m█[0m[38;2;98;153;38m█[0m[38;2;97;157;42m█[0m[38;2;105;159;44m█[0m[38;2;104;159;40m█[0m[38;2;105;157;40m█[0m[38;2;105;156;40m█[0m[38;2;110;161;41m█[0m[38;2;81;143;41m█[0m[38;2;100;158;42m█[0m[38;2;102;154;42m█[0m[38;2;96;152;39m█[0m[38;2;129;168;41m█[0m[38;2;100;152;37m█[0m[38;2;95;153;38m█[0m[38;2;100;155;37m█[0m[38;2;139;172;45m█[0m[38;2;127;162;37m█[0m[38;2;84;148;44m█[0m[38;2;124;166;43m█[0m[38;2;120;166;47m█[0m[38;2;83;147;42m█[0m[38;2;82;147;43m█[0m[38;2;79;147;40m█[0m[38;2;51;129;50m█[0m[38;2;57;133;46m█[0m[38;2;71;140;50m█[0m[38;2;69;139;42m█[0m[38;2;71;142;42m█[0m[38;2;98;151;43m█[0m[38;2;98;157;47m█[0m[38;2;71;142;50m█[0m[38;2;56;134;44m█[0m[38;2;89;149;41m█[0m[38;2;68;137;41m█[0m[38;2;60;136;49m█[0m[38;2;45;123;46m█[0m[38;2;47;128;49m█[0m[38;2;48;127;52m█[0m[38;2;48;129;53m█[0m[38;2;66;142;53m█[0m");
$display("[38;2;62;133;47m█[0m[38;2;45;120;45m█[0m[38;2;37;112;43m█[0m[38;2;34;113;48m█[0m[38;2;64;137;42m█[0m[38;2;58;132;42m█[0m[38;2;41;116;49m█[0m[38;2;41;117;54m█[0m[38;2;66;140;55m█[0m[38;2;69;141;41m█[0m[38;2;64;137;47m█[0m[38;2;46;119;42m█[0m[38;2;47;122;45m█[0m[38;2;42;117;48m█[0m[38;2;71;142;42m█[0m[38;2;74;140;40m█[0m[38;2;48;122;45m█[0m[38;2;45;119;44m█[0m[38;2;54;127;48m█[0m[38;2;84;149;43m█[0m[38;2;93;153;42m█[0m[38;2;91;153;43m█[0m[38;2;93;151;42m█[0m[38;2;91;153;37m█[0m[38;2;93;152;46m█[0m[38;2;70;138;42m█[0m[38;2;86;150;42m█[0m[38;2;95;150;36m█[0m[38;2;93;148;42m█[0m[38;2;98;151;37m█[0m[38;2;99;153;40m█[0m[38;2;103;152;36m█[0m[38;2;99;154;39m█[0m[38;2;109;155;35m█[0m[38;2;115;162;41m█[0m[38;2;101;157;38m█[0m[38;2;100;157;39m█[0m[38;2;111;160;36m█[0m[38;2;110;160;40m█[0m[38;2;106;157;39m█[0m[38;2;115;166;42m█[0m[38;2;105;159;39m█[0m[38;2;95;155;41m█[0m[38;2;94;151;41m█[0m[38;2;107;157;35m█[0m[38;2;103;154;36m█[0m[38;2;104;159;40m█[0m[38;2;102;153;34m█[0m[38;2;111;160;37m█[0m[38;2;102;155;48m█[0m[38;2;83;142;43m█[0m[38;2;95;153;43m█[0m[38;2;101;155;43m█[0m[38;2;102;156;43m█[0m[38;2;94;154;45m█[0m[38;2;92;152;41m█[0m[38;2;86;149;44m█[0m[38;2;82;142;43m█[0m[38;2;90;153;48m█[0m[38;2;86;145;37m█[0m[38;2;92;151;39m█[0m[38;2;95;153;43m█[0m[38;2;72;140;44m█[0m[38;2;87;147;42m█[0m[38;2;88;147;36m█[0m[38;2;61;128;43m█[0m[38;2;68;136;49m█[0m[38;2;86;146;35m█[0m[38;2;96;153;39m█[0m[38;2;90;149;44m█[0m[38;2;89;152;41m█[0m[38;2;105;156;40m█[0m[38;2;133;172;46m█[0m[38;2;80;144;38m█[0m[38;2;101;151;38m█[0m[38;2;120;165;45m█[0m[38;2;74;142;53m█[0m[38;2;103;152;37m█[0m[38;2;58;131;38m█[0m[38;2;59;134;39m█[0m[38;2;69;143;52m█[0m[38;2;66;138;45m█[0m[38;2;60;132;45m█[0m[38;2;49;125;42m█[0m[38;2;40;117;49m█[0m[38;2;42;121;49m█[0m[38;2;50;128;43m█[0m[38;2;63;137;43m█[0m[38;2;60;133;54m█[0m[38;2;46;124;50m█[0m[38;2;43;121;48m█[0m[38;2;55;131;45m█[0m[38;2;58;137;49m█[0m[38;2;37;117;45m█[0m[38;2;23;103;49m█[0m[38;2;30;110;53m█[0m[38;2;32;112;51m█[0m[38;2;52;130;52m█[0m[38;2;51;132;49m█[0m[38;2;47;124;52m█[0m");
$display("[38;2;48;125;52m█[0m[38;2;54;130;48m█[0m[38;2;49;127;52m█[0m[38;2;35;111;55m█[0m[38;2;35;112;53m█[0m[38;2;36;112;56m█[0m[38;2;62;138;52m█[0m[38;2;39;117;57m█[0m[38;2;43;118;58m█[0m[38;2;57;136;57m█[0m[38;2;47;126;44m█[0m[38;2;36;115;50m█[0m[38;2;40;117;53m█[0m[38;2;35;112;50m█[0m[38;2;55;130;44m█[0m[38;2;32;111;53m█[0m[38;2;40;117;52m█[0m[38;2;62;136;39m█[0m[38;2;67;140;43m█[0m[38;2;70;143;49m█[0m[38;2;48;124;44m█[0m[38;2;52;124;46m█[0m[38;2;81;146;46m█[0m[38;2;68;139;37m█[0m[38;2;80;148;43m█[0m[38;2;70;144;40m█[0m[38;2;61;129;48m█[0m[38;2;59;131;45m█[0m[38;2;81;149;44m█[0m[38;2;49;120;42m█[0m[38;2;78;146;48m█[0m[38;2;78;148;48m█[0m[38;2;87;150;38m█[0m[38;2;68;135;36m█[0m[38;2;83;145;49m█[0m[38;2;90;149;40m█[0m[38;2;85;148;41m█[0m[38;2;92;153;44m█[0m[38;2;90;148;37m█[0m[38;2;76;142;43m█[0m[38;2;80;144;41m█[0m[38;2;102;158;45m█[0m[38;2;99;157;44m█[0m[38;2;58;126;32m█[0m[38;2;54;126;44m█[0m[38;2;76;143;47m█[0m[38;2;79;143;41m█[0m[38;2;87;149;46m█[0m[38;2;54;130;54m█[0m[38;2;57;125;49m█[0m[38;2;79;147;48m█[0m[38;2;85;148;39m█[0m[38;2;81;145;41m█[0m[38;2;64;133;42m█[0m[38;2;67;138;41m█[0m[38;2;72;137;37m█[0m[38;2;74;144;44m█[0m[38;2;80;144;45m█[0m[38;2;79;144;45m█[0m[38;2;78;145;42m█[0m[38;2;91;151;42m█[0m[38;2;70;141;54m█[0m[38;2;80;144;38m█[0m[38;2;60;129;44m█[0m[38;2;45;119;43m█[0m[38;2;53;127;51m█[0m[38;2;84;149;47m█[0m[38;2;86;150;45m█[0m[38;2;74;143;45m█[0m[38;2;73;141;42m█[0m[38;2;75;141;41m█[0m[38;2;67;135;38m█[0m[38;2;85;145;39m█[0m[38;2;93;152;43m█[0m[38;2;83;147;39m█[0m[38;2;76;144;46m█[0m[38;2;70;141;49m█[0m[38;2;66;137;42m█[0m[38;2;61;134;44m█[0m[38;2;60;135;47m█[0m[38;2;57;132;45m█[0m[38;2;52;130;46m█[0m[38;2;58;133;52m█[0m[38;2;45;124;50m█[0m[38;2;30;109;47m█[0m[38;2;32;111;54m█[0m[38;2;39;123;45m█[0m[38;2;43;127;54m█[0m[38;2;29;114;52m█[0m[38;2;40;121;56m█[0m[38;2;63;139;50m█[0m[38;2;60;140;58m█[0m[38;2;37;117;58m█[0m[38;2;35;117;58m█[0m[38;2;26;113;54m█[0m[38;2;42;124;53m█[0m[38;2;46;127;50m█[0m[38;2;47;124;54m█[0m[38;2;37;117;53m█[0m[38;2;36;115;50m█[0m");
$display("[38;2;41;121;53m█[0m[38;2;27;109;52m█[0m[38;2;42;120;51m█[0m[38;2;55;133;51m█[0m[38;2;30;107;52m█[0m[38;2;34;111;52m█[0m[38;2;29;109;51m█[0m[38;2;43;121;43m█[0m[38;2;41;119;63m█[0m[38;2;30;109;54m█[0m[38;2;54;134;57m█[0m[38;2;33;115;59m█[0m[38;2;32;111;60m█[0m[38;2;48;127;50m█[0m[38;2;30;112;51m█[0m[38;2;30;109;52m█[0m[38;2;44;128;55m█[0m[38;2;61;135;52m█[0m[38;2;30;111;48m█[0m[38;2;35;112;51m█[0m[38;2;34;113;52m█[0m[38;2;57;133;47m█[0m[38;2;70;141;53m█[0m[38;2;60;134;44m█[0m[38;2;66;140;49m█[0m[38;2;58;130;46m█[0m[38;2;57;130;47m█[0m[38;2;60;131;48m█[0m[38;2;60;129;47m█[0m[38;2;55;130;50m█[0m[38;2;50;124;50m█[0m[38;2;64;135;50m█[0m[38;2;59;134;51m█[0m[38;2;52;127;46m█[0m[38;2;73;140;45m█[0m[38;2;76;143;45m█[0m[38;2;64;133;43m█[0m[38;2;68;137;48m█[0m[38;2;64;133;44m█[0m[38;2;56;129;41m█[0m[38;2;53;127;43m█[0m[38;2;47;124;48m█[0m[38;2;49;128;47m█[0m[38;2;75;144;50m█[0m[38;2;52;127;48m█[0m[38;2;43;121;51m█[0m[38;2;67;141;43m█[0m[38;2;62;133;48m█[0m[38;2;44;121;50m█[0m[38;2;45;123;54m█[0m[38;2;58;131;37m█[0m[38;2;53;127;51m█[0m[38;2;50;127;52m█[0m[38;2;46;123;46m█[0m[38;2;56;130;45m█[0m[38;2;70;146;52m█[0m[38;2;61;133;47m█[0m[38;2;55;130;49m█[0m[38;2;53;129;44m█[0m[38;2;68;139;50m█[0m[38;2;56;133;52m█[0m[38;2;52;127;49m█[0m[38;2;49;125;50m█[0m[38;2;43;121;50m█[0m[38;2;53;130;54m█[0m[38;2;69;137;41m█[0m[38;2;65;137;45m█[0m[38;2;55;129;56m█[0m[38;2;49;123;47m█[0m[38;2;68;136;43m█[0m[38;2;57;130;41m█[0m[38;2;58;132;48m█[0m[38;2;51;128;44m█[0m[38;2;58;135;48m█[0m[38;2;58;131;50m█[0m[38;2;56;134;48m█[0m[38;2;51;128;49m█[0m[38;2;52;129;50m█[0m[38;2;60;139;53m█[0m[38;2;49;127;50m█[0m[38;2;45;123;48m█[0m[38;2;41;121;50m█[0m[38;2;29;111;48m█[0m[38;2;45;127;52m█[0m[38;2;28;110;50m█[0m[38;2;32;114;61m█[0m[38;2;29;110;53m█[0m[38;2;24;113;52m█[0m[38;2;26;113;54m█[0m[38;2;43;125;50m█[0m[38;2;23;106;52m█[0m[38;2;24;108;57m█[0m[38;2;25;107;55m█[0m[38;2;24;109;56m█[0m[38;2;38;122;51m█[0m[38;2;36;120;60m█[0m[38;2;22;104;51m█[0m[38;2;34;113;54m█[0m[38;2;41;121;56m█[0m[38;2;43;125;54m█[0m");
$display("[38;2;47;125;58m█[0m[38;2;38;119;55m█[0m[38;2;26;106;51m█[0m[38;2;33;111;57m█[0m[38;2;47;127;57m█[0m[38;2;30;110;56m█[0m[38;2;26;104;54m█[0m[38;2;28;108;53m█[0m[38;2;31;115;58m█[0m[38;2;25;108;55m█[0m[38;2;27;108;57m█[0m[38;2;18;100;48m█[0m[38;2;22;102;56m█[0m[38;2;29;111;55m█[0m[38;2;24;103;50m█[0m[38;2;24;107;51m█[0m[38;2;45;126;50m█[0m[38;2;43;124;62m█[0m[38;2;26;108;52m█[0m[38;2;33;114;58m█[0m[38;2;48;127;54m█[0m[38;2;29;109;49m█[0m[38;2;38;120;59m█[0m[38;2;45;123;44m█[0m[38;2;50;129;52m█[0m[38;2;41;119;49m█[0m[38;2;46;123;53m█[0m[38;2;54;130;48m█[0m[38;2;51;127;48m█[0m[38;2;45;124;49m█[0m[38;2;43;120;46m█[0m[38;2;46;120;48m█[0m[38;2;50;123;51m█[0m[38;2;63;133;50m█[0m[38;2;49;125;49m█[0m[38;2;51;126;48m█[0m[38;2;49;123;42m█[0m[38;2;65;136;47m█[0m[38;2;52;128;51m█[0m[38;2;55;131;49m█[0m[38;2;59;134;49m█[0m[38;2;56;130;45m█[0m[38;2;37;117;51m█[0m[38;2;39;118;55m█[0m[38;2;52;126;44m█[0m[38;2;41;121;59m█[0m[38;2;36;111;48m█[0m[38;2;38;117;55m█[0m[38;2;36;114;51m█[0m[38;2;55;129;55m█[0m[38;2;39;116;53m█[0m[38;2;45;124;52m█[0m[38;2;53;130;54m█[0m[38;2;46;125;54m█[0m[38;2;43;122;49m█[0m[38;2;39;117;51m█[0m[38;2;44;121;54m█[0m[38;2;49;126;48m█[0m[38;2;54;129;48m█[0m[38;2;45;124;45m█[0m[38;2;43;121;53m█[0m[38;2;40;117;47m█[0m[38;2;40;117;51m█[0m[38;2;43;119;51m█[0m[38;2;56;132;49m█[0m[38;2;48;125;52m█[0m[38;2;50;126;55m█[0m[38;2;56;130;57m█[0m[38;2;58;132;40m█[0m[38;2;51;125;48m█[0m[38;2;42;121;48m█[0m[38;2;47;127;55m█[0m[38;2;50;127;52m█[0m[38;2;41;119;43m█[0m[38;2;53;126;48m█[0m[38;2;41;121;51m█[0m[38;2;42;120;53m█[0m[38;2;48;127;57m█[0m[38;2;35;115;52m█[0m[38;2;31;115;54m█[0m[38;2;35;118;59m█[0m[38;2;37;119;55m█[0m[38;2;29;112;54m█[0m[38;2;23;104;55m█[0m[38;2;36;123;56m█[0m[38;2;24;107;57m█[0m[38;2;24;108;61m█[0m[38;2;26;108;58m█[0m[38;2;33;116;54m█[0m[38;2;25;107;61m█[0m[38;2;20;103;55m█[0m[38;2;26;112;61m█[0m[38;2;18;103;50m█[0m[38;2;24;105;54m█[0m[38;2;19;105;55m█[0m[38;2;27;108;58m█[0m[38;2;40;123;58m█[0m[38;2;36;116;57m█[0m[38;2;34;115;50m█[0m[38;2;45;126;53m█[0m");
$display("[38;2;37;115;55m█[0m[38;2;42;117;60m█[0m[38;2;28;111;57m█[0m[38;2;27;108;59m█[0m[38;2;21;106;52m█[0m[38;2;27;111;55m█[0m[38;2;21;99;51m█[0m[38;2;23;104;57m█[0m[38;2;23;100;51m█[0m[38;2;34;112;57m█[0m[38;2;22;103;51m█[0m[38;2;21;107;53m█[0m[38;2;29;107;61m█[0m[38;2;23;106;54m█[0m[38;2;29;110;53m█[0m[38;2;35;118;58m█[0m[38;2;31;113;59m█[0m[38;2;20;100;50m█[0m[38;2;30;114;53m█[0m[38;2;34;118;59m█[0m[38;2;33;114;60m█[0m[38;2;25;105;52m█[0m[38;2;43;123;57m█[0m[38;2;44;127;51m█[0m[38;2;36;115;48m█[0m[38;2;36;112;49m█[0m[38;2;41;120;54m█[0m[38;2;58;134;53m█[0m[38;2;47;126;53m█[0m[38;2;49;123;51m█[0m[38;2;44;125;43m█[0m[38;2;56;131;56m█[0m[38;2;48;127;50m█[0m[38;2;53;128;49m█[0m[38;2;47;121;48m█[0m[38;2;48;120;49m█[0m[38;2;60;133;54m█[0m[38;2;53;128;53m█[0m[38;2;51;128;51m█[0m[38;2;50;123;50m█[0m[38;2;37;114;52m█[0m[38;2;40;120;53m█[0m[38;2;39;116;49m█[0m[38;2;39;118;54m█[0m[38;2;34;113;50m█[0m[38;2;37;119;58m█[0m[38;2;49;130;63m█[0m[38;2;32;111;54m█[0m[38;2;38;115;46m█[0m[38;2;42;125;55m█[0m[38;2;46;124;56m█[0m[38;2;42;123;54m█[0m[38;2;41;123;54m█[0m[38;2;50;125;58m█[0m[38;2;43;122;50m█[0m[38;2;48;125;52m█[0m[38;2;44;125;52m█[0m[38;2;40;119;50m█[0m[38;2;43;119;54m█[0m[38;2;42;123;55m█[0m[38;2;45;123;52m█[0m[38;2;48;125;62m█[0m[38;2;45;121;50m█[0m[38;2;43;123;53m█[0m[38;2;40;118;49m█[0m[38;2;41;120;56m█[0m[38;2;40;121;55m█[0m[38;2;44;126;57m█[0m[38;2;39;117;48m█[0m[38;2;35;117;53m█[0m[38;2;48;129;57m█[0m[38;2;39;119;54m█[0m[38;2;41;122;56m█[0m[38;2;39;117;55m█[0m[38;2;42;123;50m█[0m[38;2;39;116;47m█[0m[38;2;38;120;53m█[0m[38;2;30;111;50m█[0m[38;2;37;115;54m█[0m[38;2;38;122;58m█[0m[38;2;33;116;60m█[0m[38;2;24;108;51m█[0m[38;2;26;110;59m█[0m[38;2;40;123;69m█[0m[38;2;24;108;60m█[0m[38;2;23;104;57m█[0m[38;2;21;107;54m█[0m[38;2;25;108;52m█[0m[38;2;23;109;56m█[0m[38;2;26;114;65m█[0m[38;2;20;101;53m█[0m[38;2;23;107;56m█[0m[38;2;28;110;60m█[0m[38;2;24;111;61m█[0m[38;2;25;110;59m█[0m[38;2;33;115;60m█[0m[38;2;24;108;55m█[0m[38;2;32;112;56m█[0m[38;2;35;118;55m█[0m[38;2;34;112;53m█[0m");
$display("[38;2;34;114;51m█[0m[38;2;40;117;54m█[0m[38;2;34;113;55m█[0m[38;2;31;111;59m█[0m[38;2;27;109;57m█[0m[38;2;28;110;58m█[0m[38;2;22;100;55m█[0m[38;2;24;109;58m█[0m[38;2;20;101;52m█[0m[38;2;21;104;56m█[0m[38;2;22;104;53m█[0m[38;2;21;104;53m█[0m[38;2;25;104;55m█[0m[38;2;27;108;59m█[0m[38;2;25;106;56m█[0m[38;2;23;105;53m█[0m[38;2;25;107;55m█[0m[38;2;33;111;57m█[0m[38;2;34;118;62m█[0m[38;2;29;110;57m█[0m[38;2;26;106;56m█[0m[38;2;44;124;66m█[0m[38;2;31;113;56m█[0m[38;2;27;109;54m█[0m[38;2;35;117;54m█[0m[38;2;37;118;53m█[0m[38;2;45;121;56m█[0m[38;2;37;114;51m█[0m[38;2;43;121;55m█[0m[38;2;40;114;53m█[0m[38;2;42;121;50m█[0m[38;2;48;123;49m█[0m[38;2;47;123;51m█[0m[38;2;45;122;47m█[0m[38;2;54;128;52m█[0m[38;2;50;123;51m█[0m[38;2;54;129;53m█[0m[38;2;58;133;57m█[0m[38;2;49;122;44m█[0m[38;2;47;122;48m█[0m[38;2;49;123;53m█[0m[38;2;46;122;51m█[0m[38;2;39;117;50m█[0m[38;2;39;118;50m█[0m[38;2;46;122;54m█[0m[38;2;45;121;53m█[0m[38;2;39;118;54m█[0m[38;2;39;116;53m█[0m[38;2;42;120;52m█[0m[38;2;41;121;58m█[0m[38;2;40;117;50m█[0m[38;2;43;122;53m█[0m[38;2;45;121;52m█[0m[38;2;41;118;51m█[0m[38;2;42;120;56m█[0m[38;2;47;122;55m█[0m[38;2;47;125;57m█[0m[38;2;44;122;57m█[0m[38;2;44;120;53m█[0m[38;2;40;119;55m█[0m[38;2;47;125;60m█[0m[38;2;40;118;54m██[0m[38;2;43;122;56m█[0m[38;2;35;118;48m█[0m[38;2;41;121;56m█[0m[38;2;50;133;68m█[0m[38;2;39;118;59m█[0m[38;2;37;116;54m█[0m[38;2;34;111;53m█[0m[38;2;32;113;53m█[0m[38;2;31;114;54m█[0m[38;2;41;121;54m█[0m[38;2;40;122;55m█[0m[38;2;38;121;58m█[0m[38;2;34;116;53m█[0m[38;2;35;114;53m█[0m[38;2;33;116;50m█[0m[38;2;32;112;50m█[0m[38;2;34;116;62m█[0m[38;2;36;116;63m█[0m[38;2;27;111;58m█[0m[38;2;35;118;60m█[0m[38;2;24;109;54m█[0m[38;2;25;109;59m█[0m[38;2;26;107;59m█[0m[38;2;21;104;58m█[0m[38;2;22;106;57m█[0m[38;2;26;110;58m█[0m[38;2;29;112;60m█[0m[38;2;30;115;63m█[0m[38;2;27;114;57m█[0m[38;2;22;106;55m█[0m[38;2;20;105;53m█[0m[38;2;25;107;57m█[0m[38;2;22;106;53m█[0m[38;2;31;110;59m█[0m[38;2;37;118;59m█[0m[38;2;29;110;47m█[0m[38;2;37;114;54m█[0m");
    
    $display("\n");
    $display("                   \033[32m\033[5m █████ █████ █████ █████ █████ █████ █████ \033[0m");
    $display("                   \033[32m\033[5m █     █   █ █   █ █   █ █     █       █ \033[0m");
    $display("                   \033[32m\033[5m █     █   █ █████ █████ █████ █       █  \033[0m");
    $display("                   \033[32m\033[5m █     █   █ █  █  █  █  █     █       █  \033[0m");
    $display("                   \033[32m\033[5m █████ █████ █   █ █   █ █████ █████   █  \033[0m");
    $display("\n");
    
    
    
    
    $display("        -------------------------------------------------------------------               ");
    $display("                          --                        --               ");
    $display("                          --  Congratulations !!    --               ");
    $display("                          --                        --               ");
    $display("                          --   \033[0;32mSimulation PASS!!\033[m    --");
    $display("                          --                        --               ");
    $display("        -------------------------------------------------------------------               ");
    
end endtask





task display_pass_gradient;
    input integer patcount;

    integer i, indent, wave_index;
    integer green[0:15];
    reg [8*22:1] msg;
    reg [8*8:1] num_str;
    reg [7:0] ch;
    integer wave_pattern[0:79];

    real pi;

begin
    // 16-step green color palette (ANSI 256-color codes)
    green[0]  =  22; green[1]  =  28; green[2]  =  34; green[3]  =  40;
    green[4]  =  46; green[5]  =  82; green[6]  =  118; green[7]  = 154;
    green[8]  =  190; green[9]  =  156; green[10] =  120; green[11] =  84;
    green[12] =  48; green[13] =  42; green[14] =  34; green[15] =  28;

    // Generate circular wave pattern using sine function
    pi = 3.1415926;
    for (i = 0; i < 80; i = i + 1)
        wave_pattern[i] = 15 + $rtoi(15.0 * $sin(8.0 * pi * i / 80.0));

    wave_index = patcount % 80;
    indent = wave_pattern[wave_index];

    msg = "Pass Pattern NO. ";
    $sformat(num_str, "%0d", patcount);
    
    // Apply indent (horizontal shift)
    for (i = 0; i < indent; i = i + 1)
        $write(" ");

    // Print "Pass Pattern NO. " with gradient coloring
    for (i = 0; i < 17; i = i + 1) begin
        ch = msg[8*(17 - i) -: 8];
        $write("\033[38;5;%0dm%c", green[i % 16], ch);
    end

    // Print pattern number with continuing gradient
    for (i = 0; i < 8; i = i + 1) begin
        ch = num_str[8*(8 - i) -: 8];
        if (ch != 8'd0)
            $write("\033[38;5;%0dm%c", green[(i + 17) % 16], ch);
    end

    // Reset color and move to next line
    $display("\033[0m");
end endtask




endmodule

