`ifdef RTL
`define CYCLE_TIME 20.0
	`define RTL_GATE
`elsif GATE
`define CYCLE_TIME 20.0
	`define RTL_GATE
`elsif CHIP
`define CYCLE_TIME 20.0
    `define CHIP_POST 
`elsif POST
`define CYCLE_TIME 20.0
    `define CHIP_POST 
`endif

`define CYCLE_TIME_DATA 31.7

`ifdef FUNC
`define PAT_NUM 2048
`define MAX_WAIT_READY_CYCLE 2000
`endif
`ifdef PERF
`define PAT_NUM 2048
`define MAX_WAIT_READY_CYCLE 100000
`endif


`include "../00_TESTBED/MEM_MAP_define.v"
`include "../00_TESTBED/pseudo_DRAM_data.v"
`include "../00_TESTBED/pseudo_DRAM_inst.v"

module PATTERN(
    			clk,
			  rst_n,
		   IO_stall,


         awid_s_inf,
       awaddr_s_inf,
       awsize_s_inf,
      awburst_s_inf,
        awlen_s_inf,
      awvalid_s_inf,
      awready_s_inf,
                    
        wdata_s_inf,
        wlast_s_inf,
       wvalid_s_inf,
       wready_s_inf,
                    
          bid_s_inf,
        bresp_s_inf,
       bvalid_s_inf,
       bready_s_inf,
                    
         arid_s_inf,
       araddr_s_inf,
        arlen_s_inf,
       arsize_s_inf,
      arburst_s_inf,
      arvalid_s_inf,
                    
      arready_s_inf, 
          rid_s_inf,
        rdata_s_inf,
        rresp_s_inf,
        rlast_s_inf,
       rvalid_s_inf,
       rready_s_inf 
    );


`protected
=cL;LW)8G2XZ6aadc+/)IK;KT7JTdURFXL1CdBd:/:[F;g9#D07-7)U5;DY<WE<N
GP9ZeULAPRACXHXV@IOBa^JJO/;&be/IL[EKZf@,6cLBfD&EV?WSUA_#Y671[YKK
B-L96@M(b/G?M8LMZ_[/Ua0#T5BS_-RV,a.@MLe8JVLUa_XFIX<UIM<K&=\=OF-;
MHK.9=(d?&B#59cX4X@5+-(<N[S9/a7^dR1UU\354@a3g3EMF6cCdOEDO?FI;f-^
9YCZ</T&DWb\6FK5_LKg+;;)7?QJcecII,M;>K=I.MCB/]HA&c=PC]UJWF8YUU73
aD(4[N^eWYP5SN,XMN);f/g9ZD+PGTdR)V0cO0M)\^4B&@K-=8dP8ZB4VG+H1fR1
SVCF3dXD0>RZ/#;K5S\#L&-G\ZX<?d2+@$
`endprotected
output reg			  clk,rst_n;
input				IO_stall;


`protected
?b;D.BZIdP6cZI7^aZG8UYfE@JT;6^3(H&PX^>,,(d__Xa9JBK]J))>#&N1?Z]a=
CK?e/BK&,+N0Cgg2W2V3HaGe5O]296>a^[aTW7??#=X_G$
`endprotected
input wire [WRIT_NUMBER * ID_WIDTH-1:0]        awid_s_inf;
input wire [WRIT_NUMBER * ADDR_WIDTH-1:0]    awaddr_s_inf;
input wire [WRIT_NUMBER * 3 -1:0]            awsize_s_inf;
input wire [WRIT_NUMBER * 2 -1:0]           awburst_s_inf;
input wire [WRIT_NUMBER * 7 -1:0]             awlen_s_inf;
input wire [WRIT_NUMBER-1:0]                awvalid_s_inf;
output wire [WRIT_NUMBER-1:0]               awready_s_inf;

`protected
P-XXY^27\dd\1;P#6>KbDdOP3[DDKC4YS;Ya&RNZ5gB_;;[C=\/>.)9@W^Nc?YKJ
O8VUZTa+095YOTE(d_^Wc)TC\O&6FbLdUVdYBF3ae=I_D$
`endprotected
input wire [WRIT_NUMBER * DATA_WIDTH-1:0]     wdata_s_inf;
input wire [WRIT_NUMBER-1:0]                  wlast_s_inf;
input wire [WRIT_NUMBER-1:0]                 wvalid_s_inf;
output wire [WRIT_NUMBER-1:0]                wready_s_inf;

`protected
eO-Ha61<^=9bGHSGI:R@BGPZ;e\XGUZ(J,QO8gB2bII;^-+7[QcN/)SbL&dLEAC4
@]<;U8QXeU>b</:&a0Z/>><-3+=J5GU22ZV=MDP>2R^;G$
`endprotected
output wire [WRIT_NUMBER * ID_WIDTH-1:0]         bid_s_inf;
output wire [WRIT_NUMBER * 2 -1:0]             bresp_s_inf;
output wire [WRIT_NUMBER-1:0]             	  bvalid_s_inf;
input wire [WRIT_NUMBER-1:0]                  bready_s_inf;

`protected
H4FF=.>8NVYA^J.[cSNLJ0.3f<U>ZK8)CE9e-)RA<5,bU^,Z>68\&)6(.2#NZV)S
><=cedC(6NPBD^@Ud,LV#fOCOS+P3X[;TN^?OH9UL-eWXGJ\W8J).NI46g8EP&1O
PMf)+I+<+J?;W.9)@VP+#LOC8$
`endprotected
input wire [DRAM_NUMBER * ID_WIDTH-1:0]       arid_s_inf;
input wire [DRAM_NUMBER * ADDR_WIDTH-1:0]   araddr_s_inf;
input wire [DRAM_NUMBER * 7 -1:0]            arlen_s_inf;
input wire [DRAM_NUMBER * 3 -1:0]           arsize_s_inf;
input wire [DRAM_NUMBER * 2 -1:0]          arburst_s_inf;
input wire [DRAM_NUMBER-1:0]               arvalid_s_inf;
output wire [DRAM_NUMBER-1:0]              arready_s_inf;

`protected
eA8AA/YQfX^aP4>K<LK@R;W/..TZ4g&g6g4_ZLb#U7f>8Ec==.YT/)AX+Sd:F&6)
YM.O14?T=.2aT+R=5M=/A4ZT;\S?&3=AF9T@E6\P_U9NZU\8?3:,]]If^U18@(;9
/C/;G063,,_Q_1>ZC/4AASZT5$
`endprotected
output wire [DRAM_NUMBER * ID_WIDTH-1:0]         rid_s_inf;
output wire [DRAM_NUMBER * DATA_WIDTH-1:0]     rdata_s_inf;
output wire [DRAM_NUMBER * 2 -1:0]             rresp_s_inf;
output wire [DRAM_NUMBER-1:0]                  rlast_s_inf;
output wire [DRAM_NUMBER-1:0]                 rvalid_s_inf;
input wire [DRAM_NUMBER-1:0]                  rready_s_inf;

`protected
2&H<RO7&3_)c@Y]]UP+NN]SMAbbZ_<+3>,V/)?X>2@?C+g8&I[&+))E)fL-,E2aW
>:FgO6a+./9[O5I+<67.:Y:5LQ(UPG1eUQ\5UdXYF\6e.PGc2;50<:+;DDN9QK58
)QR,D^A>;a9MI)=#F?3OZ46aaT>+@dF)8^&deE\<OQc3fNd.+LbD6)7)VE2@H@;2
IN0]d=L.\/5+B<dU=&W>KF/gOTI,._N+K<4\]7:8@\<.U8B,d+CLM2PBa^4dRGP,
G(N+Q7)NOagf9CT.#UG9V>6@UY+O:Te.5a_[RH4CG7\XgC:F+V#/I>C?ILKZ]A7_
N.K[5PKF=UZf[:)>;Ng2W14P(>(SYP1bdM;6APe?7MX>VINHPM:DCXW=@8C_<U>O
dVZA_U?e-D-W+2VIJ+(cG:.\eE\J\8T,V^P93XI7.I@c9+4IbSZ#/8M?1-CePG/,
Y<5ebW84.)aTdY#DD/PQ(S>?-^TZOFXC9b0TV.3_[KY&_CY(2#X)#]0NfNB&Nc1_
Af9/AYLN?-?gN-XPD^<1Q:\=><E[O\AVXaf,a,Z#+23#;&fE46]4^.4L2Td7adab
T4P65)A?SPdPG#1[eD6KcGT[PK-+X@5<IH=CAf\>F=eRSe_f.T]^NE?OZgZ9E&MS
PdSPM8_cCXVQNQDQ>W5c1R1Y:VR-0_/5C4MWB5_D2@>dCRb>&0c.bB7]MM0P>/MC
22U42W=5>,;fDLZRA:5b]5DMgBg=8,U(c8V:a,4+;+,<;]0#KZ#96U3P-/[[=FD:
53VO?f62>)aFfb.4M.U/?NJ&WURBcRWD=,?6@R3cb]@bDdPF[a\F2PJ7XRLY@c/>
NgdY-O/4.KM0aJSV_C+ag5V?CAST7A@GMI.LCY6?51fC5E81RTC)fd@_4[g&,F;c
K2.DHRL?@)QQF^6<[6Q.QF]/.;-PgT+BC/ZW;[^0V1KYQ?bbQ+.S4^@BGHYedYVC
?76+=UDbCef7>07I5GOH,-3M=)(,Pb_3>Q-F6BZaGbfXO6IK4&1->X8@TD9_2O+9
?Hd(A2c2dE]DaSg\SHH&CbMS\BE.(-XgVBIHMS0,^&KUY?L_TLMIc2\Ed+QT@LRB
Y=,D?8<--gV>N-;==FRGGAc?_>MA[&J-gJ)X<;JIPE4;74UIa;&H=D3/)f1)g&R=
DC_^F/Sa]Z(L-2,]]B:Q8/>JZ_X<;f?H]:\I&H#,,=]\Y6B[^^)/JX3@R+-dTN0M
J9A2H([d/-=:ZDDYI<c/Rf9]TgWVXRb71M,a2<LTHH&T6SL2T8g<8A9YEeFE73>P
D.\5_#WUbT+\<A_,-b7\AY<G0D4bJeP=W1A?0^dM^P]^//7N>#Z.4aAZ@c1F>@.7
.<;<:QA\52O0N-H]\&]58e@I,>eO16+E^\->S5<D<7Qb[:;643<]:[,1aBLARcgZ
4]V\53VQ\]MLJAU@+b<Y-8X8/NMRb7;3D;R&)5gY@.@^#^HKG2Nc:Mc600DNc,M5
U7GIKKAC9LNLQMfgTD,ON<P\6G2-D9K4O_C#M4X@_R--D2B:K89#GL+S(gT^3#Ef
Qd1T;PEAB&,<+5DZg3W/X07(#/GTJ0=N=X9L8(99bGG8&/S6A^LALSNa>@KMJ1)X
<T_EYDI<AgK+f(cfL/:RR[-JN,8B:SHD]I]dM4>WXRXV^\83^Z-:79N^<K3_^I5[
U(@-+<WEJKCOWfK\<YUdaa7?d7OT1L)/fY\#^4]T5;gRCB,C(c2>@EXF;=@-[B-b
WLEb?G>NH1YfJ_84PY?\NDc+6cgTDTY0(O5fG/STI]/;5[:RVcH;fHa_N^&bQK-Z
dQP>e.=JCE]5G(3\dQ&09YV]IX@;B/L?c..GZ4MV=HD3_/Z<U?HVU;M/R;T)bf#<
W([>KegU,-_7f,V1U/>>Obc\ecPI^,4QO;1b@cd4HXc8OC(FUB(X]7ZW@E@R-f./
TG8IP>F1U0.&]8E9bPda#,NY<^MZJ#g2Hg+H-OER++M]7(JM<<dM#dCNKLP8AL9?
BT>(#6Y/W^&],6BeW6^)R-1M)ZN+dR#W.;[J:)FO-(LfO6^G_P+1;EgFZ,aH3G-^
FL/bbCK\#9KdQ>QDR4DfVAcC+S\7\F2AGO(F[YT5RCQ,<0@>WD;g#?c>KN;PK>+B
O.31??KC>=CVHLYK;-5)B[Y;SB&6B3R^d\<fADHB?[H<X=d&d5<N/Vd>TIGMQ3#M
BBePP0FZ1YTPZK2>UN<&TE>#0^=RE(If+WCcc58cN@(3.+8XLB+9[G=Z)--#OWFI
@FV@gb-LP-2J+b\T44QW3XUZ93S#5_B?X3IZTacgMK#@F5\NBe?:NNQ-CFL/Za8U
E4J_./>J2eST.ZD)9QV[>K1NW#DAN5]]WOa4\.A1Q.B@T)/]bZ),I415;a;?Q/.;
8\Bb[&K)MA<<03@.f0Fd29R36IfD/N,90FTg]^/KU0,FJKKdT(J+g2T=SXCUge)@
9U/AJ82IeRB47M\[KM/WdaO>J#1/5<aV1gK2>5dY;1UPHF;@5c^14a0Z8K&@:d0#
WW78VJI)I><^O;[RR-<RAMN^7cRR+<B07@CbKK+D5(=1fGdCK9[?8CWQ]X8L0;0+
;e=IVLXL0/8>3L+US:W>=R2_J^F.90CU+GKOY+TA]1NOUT-\Q#[F9L/(:CG9d?I/
;(1B.EL.B]-=02(U;]a+[]2/NdXB+1SPO&Lg2XP+/)6:37:ebGUJ@L7Q3GUK+BT:
QQ&]X&H3@LO0V9eHf)EIH(I#KU0-.XD\GV;C+Y,C:4d2X2dWE;(+cK><<\/8<8U@
5RWKa])A[B3JCG434G=TS^3HTTY^a7/@Nf2b^EbY<Z-Bf,DTFB_L9Qf42M_K,<D^
.,Mc;AE_M?M,G&OJ<RJ@=HF/&-(R]bM)MC]^>+XgTTT8/>B;bc8c[F6c=96-)8.E
9FS^e@cV)CWP(95c&PbAVX]R[?]MX_cS.&gWbCU6c&C5]5d1RKbUB:1BTeRH6E3+
DU[B+^HNW=-5J6f+7Y4CYJI>Pg,fTMU_[0-ZPDI95L.8HgdFK:da5bC0./7SeMHJ
<dE;P=eYUEM2D0,)LHI9BZJ#6=E2DZQaWZ5PPTUeBFBZLDTW?J;Y(Jeb\D4IZa6f
<SSJ<ENV,5d:X(Y,-AC]#Q[F@;2<(OdRA6;@dIZXP-7DVa07dYWPZS19ZA>PKKJZ
Ka<LX\^U]#U1.-C0.G]?EV\,H2-I/^Ee+e1.LIBREN9UN5^#dO(ZZ&2Z(eS8(7>g
3J3:dR>:D8T@7+5=b-dG_BCFF5,a89g-C2;K=2>R.O,,g_GFAI^5YSH<:g9O,S_,
;+=]#Bg[L/6R@,-G&=3>(bDI4GgQ^,D#BHfRg+];MLPW+6@V=29_,@XMTALD39\S
H783>^#U?(4)aca\EMc9,@RZCL6]VU:V]8MaP8G?d=]ETWQ6F.TO#RTO1A\2K+gC
/XSD->fa_(EAZ[LMR]?,-12R2826A-1-RSCH?aM8UaUD998?H,PGO/61&,QaF(I=
.T2,V8#?-YSH@BBU:R<Q0?;\JZ#3#R22@GXASAQSEM3,H((MCH>E,RCRP5M81a8[
UB5J(g^PZf-AQA@&X9R6M:-KNSEbP.&F/W:=K8,Y]Of>6I_)P)2e3]W:9dW?M#M<
+TQG]@De?(f.X1F;[1_fO>.(_K=,/I11/+bHV.Q=I9)H+Z>^AdL,AY@+C/1YH;W+
\A9;A2QQ?0(/EZ[_BMK.4Z(<5<,(f_G<MQVC9fP7&H56(8>DZ)WcLZ<e-^-JD_M^
\T>c^&)/04=S1_I/9GLH-OIO;fJQW,EFIFPHP)fNY)AN2b&,=2MecNW+ICZgSR4Z
0J18&>Y3Z,)N590<<#ZB6ATYBdb1C[QH^FQMQ6VE8c?CGadU,6^J-D1NV[7E[/dH
+FZ-[0M,R]C@^M>ZE]KfV<OGP2(EDZ@NV8:-Z)c<(O]FLRIA&-F]/Hc)(0=_XK#&
IZACEM+JT40YM_L:=VEVJ/7^,8N]BPg.R&f?YNEOD?9D.g39NJT^DG,2^3cg@TCD
]N0-g8[:,:83NC)283g_W0[WDI\?+T7:Q1\gM)9YJME3?bBZQ;B5Kf2-\[2BJ^#6
V>dX[M5CML4(\#9TVA_@-\Mc9N4f(ULVf^K2L\F_K2d82[BXWF)0cL@c)P.#QGXC
dDWM\S.ILA?N80]<8;bJTS[;Ba:5.R@=3@H/c.baOXZB7UeQB=VK3H@E[/+<>aP6
Y).VKf3@N9OBD,KL6&[#cS<a(4(+<IG=VF4-Ib:R,??Xd1e_KM--[F:<c24KTJDT
TINHAQ99W(243S8->\TL^UC?]aeY,8fQ_^LC>G,afR^_N(&/6NJF27H>[<(L_WQ+
GRU8,@1&\>\YPI&H]U\#ZaC(+XdaD3BQ0fQT]I@c?;H50[4UE4,??CY\@>T,,<]e
+6E0&e05fK)HA^V5aYf2+?=)+<0OE2/g3YFc)[C27[O)F>X>a25Q279@_<U<>_d)
^cD,E-@c2(\aX_AZG_NB6c=Ud#O1G.6_IcX,)/Q&-]AX98+)P/Ka8VW.6J=UJQXP
Z)7R&M>G:e92Bfb.c^1+Z8<H&gJHfQ++A82WMIY(7\R>Zd76ST<9DA[RGWXCN4\1
1DbWL7@L:.\VYG3OH=f3f=N=@#RR5R60g:XTN/VXTG+,f?W(U>(U81I\U)JDQN&_
EV/#ML=a2_U]QI/N08(PHC]I-&/55VbO1W(b/FYa[FDg^HVT.[cUFQ6aBDU:[0CO
1=gQ+2+K9?0W;PZ>N<I2GX=Ed)V8fQ@[TTE+-J5D:?^V+&1G/-[A4IW2277Y=SXF
NcHKIf[B(;2;J:?>b<^9(eW96cUNfXAP&,_8KZ8ET(@:C(&-P/EPB46MM3L4Xc@:
c.V=KZ1b2-bL8<PXER7;gfCd97[YJ4C5&>7aY^5@>H+d:97=-]Y8NH/2dcIgLX-9
^,2RI]bbG:F\J-6/VUXX;?ML4R.f==&Ta-K0UR4SE:[/8ISDJ?b#c<1_@M/XWVV+
UMccAUD?9EQ[^>fAM.\Sg;^;&IOc1Q/=,FX294;H^L=77[+=/7[&P;RG@0H2cNU[
N556)H:S_ZfNdLg4g^MX^:Z#ZY;2\&;5^Y;W]N./=-W8[a)LHUWd6aOR9\I6(K6R
XZF&,O-=_>fN##3]O]]1?^JQL&K+\\I2=(b^,Y&R^LEaX:XD,4OE8<6?aWe/W1#/
QRQ5)c<\2[B/MFYQLJC,HfZA@V;]NY44QQRaJ8+M>ccb@a9YUW(7KBV2ee&LC(D(
NB5[=BFO>-DI4M4E-6_P/+bQ9W>(\MJHe^>@H3^<</0),Kc=YNSZ/Ub92#&<XJQG
I^Tf=g>NR/e>R6]IZ-b2W1U;M).RAPMS..2b:c??96XJOdK2c]9#fg&D29TgZ4^^
>Y5d4+@FaF\_<:5L]A3_KG_-0F,6=ZL[16cA_NG6A0-/66;DQEf@-&PecO/86R+1
E(c9Q3Z(A92/d\])&5-b(I[[@0_-QO:MPEUFXT#:(K#0?EK51_c#R^J27/dN:ZLL
.MH]6.DD;(eIT6X@4QX)0\,:g)@-#ba9H8PT9W<&8QMDNab7X2D(.41>D)da:g;A
,4X60.d4>\d.=6Q>_CG+,g&-H+I^XI@^NPY4805;??CCM]<9[4T#Z7TKPG;1V/16
@Ag906P9D+&WEY42g@[+gLQbbIVC=8#29Ae/-^J24fE>5I=9M\5][+VW@e1QeQD.
7(IHc3F]L-g(V4OK]C]VWYU>HRG3-=C@eWQ[+dJG0B#A<3=69,I;R>_:2>@MHHV1
<0SW2cNWYVQf;.VSa383(R5;)DDcWa)Z#N=#CDLH:+X(T8EI?YCNG7R_2AL8O?2<
YH)cC3\.)IJJaR5LGcad(0PUg1@Z4@#Kd\KOFOcQI>WcU?/X?=.QC4(/Tf5CW.65
V([V=7++.X+F(8^_g9cVSID>W,^3V:W/><&BE:GSb^S2PZb59I@Yf).KD+RW5KT]
BO8N#-cJ?:;/\<fQ_(36_X(LKE(\Df:PD(:3]OVN,_da_P[5gVX6cAgd53b:2fIb
DDG.B]0]GdXL/Hg@]gT9Q2Ff(V9c):JEA7g9AEW]-A2:bZU>C=P3G]aEbB9RJ5O<
D7SB<4V\S=N9.YNI.aF7)NV[H3YFCe@6A-SCBW/dc6<FH/ZQ[(LU7ZOg(S>U3X0c
0Q-d&S4818OIDf1WN[58?GZL?f:<_[U>IXGe3P8QSPUT1+3/2OL/E(OHPdX]-AHU
@;SC3=f]F\^9W00a,<&X_J?dLPJ#SeB7;I&>4(dZ;MMAbWH=(0&dGELL,IO(:L/I
/NFcUXRVZXS6\cZ;Ve)1=FS<c6PF#[E9GeBU]Q7F8b+f<Qf6)I_:cP,9G1,:QL#d
&:>C<&g^/KL;3XHL765XB8.T/2ZDfWXgf#V]6(8?B9[&JFb(KC3LSf&Z6S.9PK&:
7L];b#>c+_?5f2ZU[SWbdPgY)L;,I>fGd]NgaO[^gdOMMAAHYN[4=CF)eWde;Se/
QZ]>E8cd_RSADfDBLF[(B2F;M?D&F#,fW&e_XVC97L-+KK0H]#.,5/;Y1@Q^cN01
WWIR,A/efWL8G@c5PBGU=9NUQYf;]K5Q&Qg]^4#L\K6Wa6Z1(^VXg7J\7..0T0#J
=4W9aHQ>]G,,L.&.af>U[bc89<?CQKPGGX[QP.c[2=@d@3VSWYC_8JKVIG9S/#M[
d^CP-IaP/:+bI1+Sc2=[_5UN,D.]E4C?;+:0<e^d2[b=0ff53^TcC?R&XR+OReZ.
>AH<04?]9SJ^C44<V?>R0>^9QF;-Y1c\2g&>##V.Xc,B.I3K;9Z)G?_C<#0RY\b[
Y6[<=E67ISbdC.O7cZ1f+U^)]IZ1Z&JDeVP<b/f2::9+.6a6@,FMMX_/^004(S).
gE6/J[CPZaB8b1O)g2F7@O,-VJ\8K&<@K=b]5)&,2]dII[Jb\2bfPD4SLdF,L<_^
dKWZ9g)=[_QBPI]d0IB[BL#B/J4>/5A98GNX^+HaBUg3IYNb\Y>L?g[&B0E.7VJ2
EFLZ+2V;39RPfecSF/WaI;R/#54_YaDW2)cP[/<>?\DLefROC(Y?664XNZ^PX[A+
SUYOe2P3Q.B5?\+Y@7[f7>7J:32_ec]>@C]@=ZM]e>[9\Yb[b9fDMQ8L7P:A4>Q_
VL+Eg>)S+FX)e,E3?13T>M;IPN._?-HgB>,Z25@\3#7W<(1JMU3CS1/@QOF25STd
6Q>TR?#BfTMXH.LEO)QP]+B)I>LXgA=U>M?@J?,ZRdYY]13R5M&C&(:]VZ1b[KeJ
M;QVNKcF^H@5O,,FJ-VHZ?-R+67R;^^+\&M]0C:Bf(SR_eN283MW_fX-d_<O#&T@
.(:0G1Rd[53Q2S)<UQ;9TX+UdG764]AKa?X<Qd8f]^OQQHD/0EC9gL)HTc8<4.B1
EEUbM^?505T=3dc,?PQU(MYMY48?49]N8?O/L=^YX+YVR29Q7-IcEDR3RS_90B3_
GI2/-OOeL,@KE\1A>[LZ?H_;#V@ENQJUMf)GK:S(:NEN.>Q)A8@BB.>,;>VSd[P_
?=IfL9a<MNNJO:B-Y2CY_LU]3UX;#I_H7/O:dT/3aD\1-EL6L-^IK;SL/7Md<2?(
f[/8/d6)]&LZcc#([@I>TU?Q^.J#(MF7;JBET>4J#UZgK&f55ZFeB.Zc?fU3)7^a
c[#(4b.5+<5PgMedTM\)PY#5UG,AL1NE8O5>1AC5U??=_c-[+B#Q2a)LGJ+.&&&S
7KL9Gc1YJH^+fB)T6AKC1-SZ7OWa<D^,Fg<ZRfCC\EIdU7cQ?A+b&TX:TP6T6PIf
ge5EO@ZYX7_?6)C@?H\F#:/)8cKbc^L#LHb[.TTa6TN1H1LLA<:3\;-1.f#F71fZ
5NYfe3;fJcM0@69#IE:^1KALd#,?HZE9S8SMX;E5Ha9K_8BTED.;N+KfU[>LE>]f
=QW/CdLVFZ\^Z)CMK\\eZ;\5]>)3aS@_712)VQ=:^dMBZA/6DV_AI<,./6(-E(C9
#=cWAOH]@<aKO]2-:23JI8dK+7@7TM.Oc=Z6E0YFIA:65)Q^1Sd6W]WWU0;/J_b<
J=1VdA(&a_+^T94)AK=WN\4&?I+\aHL;Lg\B;FFI\Z[08[fLF#V^;X.KYNL&40I8
_K_/G,QP5/63NEc][<P3QT0F4G,NdDNL?[MF&<IYHN3-@,b^VJ3dEdc(/Bb;ZGUG
@?Q5bU_efS14I/7X\&\I?II6O?W\V/Uc+bR;=/\C2E.A3@3gcPEgKIEH<N/^Ie?Z
2271\HaL6&-:IMD^3TM5JGC:2<c#aW0B>1@dYd\HRRP^:-aIZHR;CffE.[MZD15[
]^(cQ-P(,<,9)WOYdM3JPO>FAXMBT)E@H1X28H-UDd1-B<ad-^.dSS8\Ngc=F:d?
HgAMWTJd2IGRcADR\Y8&WN2f./F(,bMK^M\DXA]=@0d?)C^^._L.c]SBJXRQa5>M
GQ:PL3a/aaUUU\]W\TcT65STSYbM>2dX6[M.+A-c;_)4<017U+NgT;Ja,XgGb^e,
M]^[:1_R24bVVd792D/UOB-\([[S@[8X3#1TAAGAFC1ZRDA9HYDdRW<e9)A<E&Eb
N1K(cV)eFOa\ERBaPX?C;a9)4PCTJ;&71CAUY+FEISEP,>I@UOdV6(J<(K^_dNA<
DZ7[QF&W#,[:]3?#L;E=^E@H3#A6S4=)RU.[P=4Y4B1]6?/_5De-[I^-)P[1>/>M
943>_.0:X1dGKJQ&QU2?XKdB+VeB3^fI[cIX?_QTY]>HDY=R8H_JMg:HVagGd4>H
Zd:^S.7>KbE@dNAf.GaPV@&V6,U+,fVX,)14CWU^I=.0:929AUeW,EYN(+4S1b.9
=?>3KfA?gJI:OdKJ&X^eA6ZX+IJ2UKeASW1eQ2SV(MQaUR_C@3Z/)a9[B:S-,,4\
@RfA4]-HG<FEb2E@4S8>TQ)\^:b<Ka3]2\RNQI0b-2ML^a\_.TBG1beRQ3KAWM=1
7WD^LbH?:W5JD_OOP\^-W6DJ/;5K6;J6]^:N/c==\:_J]Q(bF2+4)/)e,D26,YM#
P]>UW(Ze1A+J5cTVID7#Yc3\(Z\eeb/X810Va(NGD]7GR.2+C&9F?LAS9BXPK2[E
6BWQ[:_<(LLJQbY=/aOY]Z#[_+]2Sf(:Xgd\C0?R8E]F8E\P^MH&.0^]1UW4Y2=5
b_4J>.0:8eBeLEf3F9R-,>Zg:b>2Y9NeEgbKUAP/HXfd-1V.b[dA)#/0g1Q6,WcM
SP>c<T2BD6Ua^][7#)K9?JKY?#LLUM<N^7fa[CbG@5TI8O2:,c14EE<S\)?PH0/O
RKV<-XKERYgG<-5Fe\]/_HR_dD4:<L9<eQd(=9Z0-)fV)&<&:BId?L:McdS0\#YQ
PUXEV]:=.G/L6[M0&-ZC@U.-W[&=R3FcZBX5D\.UR.7/[6HKbbJBC4X1]\gH,H@1
;R5JV1:PLfgU>B&>B\c[KeVIFfeeH=B)XI79J>]X,(VLMa\-6XUD=X.OfZfB)#0J
DX:V9BO)#KSL4-,NWe0PC;L_,Wa:9aR&0(AQK(HQ?U#(&3^ECVS(^+RP/S;H1>-,
QegXC]5YNC1]P]XXGF?)=-20b6;I0f9MM?gEgcaZQY7P5^87NMI7b+SPJ:7\c_cA
P1CG;;H)KTT#UF:PO^Rdc0=H>^5OgNNEb->gQg.FgCAI_>N8NH?gfbT&UW[7QX&&
f@#Y1GL2+HMK/&J^Z?02J#WP]N[1\aM9:3A44F,H;8DFZ&;#]L&R:_gAG6NW;N8(
.Lb^^S)&2#RB:[_IFWYI?/QY&R&4DRY;/^AP[+[<5IT6a25CHa?].K=g[@,FTJc9
6BLD:92#,7:G3X=02D?fbD0KJ/OR0RJW>@PKEcUea4S1K75MO[^QaP>HWBB@KdET
,O^e1NdQ24_T<:&=P44ZcE)GO/OAMMd4I8ea\4?;4fbb;#-P,^4Y51;g.FQBZ3BG
b0@WVZTZ3Qd[0XT]OZcU@ZEIdg:NP).c&I\W/45_b1YL17)Ga-]+>JUaQ14PVZ+<
N\)JL.\101P;-CWHN2a?7HcR&1_OL><_ML\_#fR5[8H(gKF&e)8\DK](:0>V2?6:
)@Q[/[5[\bLD9(<,,L>VR(+8HAK_5?1AWbDUT4c:/IdW3INC#7E0Q2VbV2H0FJ-2
4U,V6cO+JSA9;a-e/-FH6EY\N]?XV]?YAR\C/@>HJ154LAX1/;30@ZZRCcdeNJ\D
R-0f#)8IO1=@T<C7,7)=T_PS4RI=7I_UZO_3K8)ZYZKR+[V+?RQ7NH4C&LM/IDVP
]UZ-.[g3+-Bf\9QB/R[ADDA&Tc:UZO02[DQ3DCB6d1LL/^::I_J1_S<GM;eX(/T,
UFe?<H2NOF)728VET.3@OG7:=Z?2)MPS@Z7?)7cO/)0DBPNS?J[97B+Y]ddA<3X/
&WT_9ILBO<b>FS^SZO^4R6Wa3Qbd^=7<UPR#+4/G^C\2[NQM&NgbKH_[8BSa]7O3
>cD+;X/Y&GG.L-IJcKKd@7:#+fKc5F7</WH8R7V^g.@TB^B?CS<d>FS4.b?EC;;Q
X(#H@.?4aDQ.D;C981M4,#S\7:/IP1JgC1-XIa#U3P=0\U@Reb@D?JFUbENGCK.-
GD(JZf80?A(OP.1,B<O6W]RdCP[I#Ld&0L;9a]d(ED)Yf>8^(UN?9bS[4S?BX1M:
b>J^[.cBIT5\<)I1F&W4Q2NdQ7UA;9/]H+5>ST^QNKPZAI62T(g&5L3I8@U1X90/
f\E.N>>HM(fb?37Ld#e+,5EWQVQ6W3=E#VK]&/&a@gE=&S@aY9XEe1GRFa#9CMeH
<SQFffdRf4PAQ<4Qe9-^MM225g&9_H@->Q+F)&cK)(6Hd6^-82#b[-R4<@Q+>3RT
0)\Y=<#XI+T:DGFdVc+0)Na_Y,[/;#_]C(?7\a\fPSJ-WB&CUI-.F^FNb9WLT5a=
HSfXfZDYf>E1M7a93,[B2YIY#.4BR+YaW(I:[2eVZ<L9HTOJ=X/5\gJc&K75ZC:<
H>^IUO/e6[FIKZ[0]0>]J+a6]WHg5W1D.(?,d)(Z5b9./D8b-\4ZRN1LW5,J=S\#
Z0@HETLea3Dg:XJ,H>9NI.UX;e3[bQL_2U11(,e.P>Q\VZH6@UJC?T0a-=;4>#K:
(<B[_,TfL)_AUWDU_)--a]>b@39a[AZH4e<4ER;6?]UVQ&3GcP1PJSSB/<]>W#Da
<0V[)]Gg-fO.V<0]R.4?978F<AP@[X5KI@YNd:0OAFc.RL4550&c3IEC?^#YZJO9
FV_CfQ/>FX<BdR3dYAC9QNTgPBX;bgfdMBXeZ:a6JdT9@Y&XY32a#d1]KP-:0aWK
WFJ4(M^&)34P7W0e^>ZZ0122;-A?a,GJU)&XFS4S<eHC&IS]_NQ-__CdfMA@MRX)
f;C@HZ77@2Acb,#Y>8d]fB/.8[>05QQ@71)AJB)L&D,OMaJ8eMgXKRC>EVdD#:OW
D#&Y3XADD#1/?93>gU#AOX>KKSgdDB(_:ZM6Ha1Gc>RA(3^P@7,L^cI:e0^_d)^=
>2??LY\S7/O-@DdYPG+Ae;a8TK;3TcCKD;=A?(_IRB^2P0@eA/bTUC)d)]--77S_
.[:,)KRK:+5YF5c=I5UV1dgbF.X3H2Vb4M0Y\MFNQU-ZW<MX4=BZ_0<)Wc\I&gIP
6&/^LF3K1K-Y_J-6F4\CS&93LJeN]&ga:ZgSLZ>7,N:>TQNW4PI3(2MJDCR41/;]
)[8]OS-:>W0.8,RVYRYC;g91\d0<6DgdZZ9Z2)>SDU0Q@2:&H[<=g)cDPK^?\5S)
0+B^A8+Q.\Z[+eG<FX?V))HFUCEY52>W[T;fb3K3aTSH6G6(Yg+f>1XA-ROC#VD9
9CV+\E2Re8TFA,.[/)/fQaU(OG>[0dBH:Y]9Z0df9.aObMCL,e^KW[3Q.+gGPY]2
Q^,+8JB0eRAa^\a@7AD7LL1VIMV[FT60<TAU#X6D(Q],:]S(+\ZF4a1_U:Ubb57;
=[e5?aJeLPa56aS@40@BE^KZd6+VC.G8]>TeV=)36cR/P]N.+E5.(E>^VKg24Xc0
M.MYDIKATGWJ_gLcQ92-#/=#R4Aa8D8gLA&[F-<caDa_^b;<+SL87L4E&<AV-Q1I
e(35Z#B>JV:>GWFTUB)H@<a3fLe;2X66N9:W;]&[UOeDPQOW4DXAY4JCAKE>,&>f
\MPIQ<A84RI[=-aU?&MAJ;c0@[a]D9R0]YX+eV5XdA[/:U7XB]NN@4a7RF#35H#V
C,AbHCYTCWf@#@BHU-@<?-M-@U-0gK2gU=Iedb-MRfS.>@1bC5WI)&UNF]&S51&,
[OHd_&dbb5>[V3aT/^MOB3f@C71\XBXR6-#aEG^IbO7/&<55Z,;5.L][3CN6+JHL
@Bf6@faJC&R-6F5,TV[<^QYT+U/L><e6eF+C]E[>9=E:c\]2CJ@CZ\Y8bC&eIg6O
gW118ALc?\8MfEC/6AB5e<ARW\B2:XKSSON@P[^P(4)\g@d5AWABGYaAK)DBC.3E
BC7[S&5C@MXSDNE&(Ig1Lc;aC;YD6VJ<N=g98=FYLESI8Kc&/[c9NC\Y5XcB^@/]
;^dP<[U,e5XWV(Y^.MD&-_>@>>MJ\QCN@IbcTCJ:0OTaI,K1VT2d@5K9+aG>XR21
?/D:940VDg?M-]QBZa1B[FP\XO/aIfTX0,6I1]1<1T4)UE)ZX2dB=->SSKOJM/09
H\D.5];1N/_d1Z[e7PA0)cQ)0_bN,;21XG6=+VO_fbZ>LegUCQF.^B[11]?2UGFc
ZY@PF7;,CM+DbM0XTb#.TS&7[)_.NeL->BAfP<&.Ac#,6gO#X9^I)Da@,J3cM1(E
HP+;Af_BRHVb?BARK3Q[]QC4deN^DY,O?0K=YGWF)8[+#)P0KF^T)OYb5,_4F](V
G=)]19EK<eN1TCX+N:L9RP,34\2Bbf&1S.F^-eQ,TQ&[L]/^=gLb>TG)6F1X?e:(
:S/L8CYEbG<SQO[ggaN,@IJK7FEVW.XHSR1?4F-HBH7]BZ?g/005bC(J]O,d5eUI
#LZSEPK)<0JJMG.?V3P?;JYR\7?,5FY)I?3DBf<3K8P(G4EUaGWXV9c=J><@/@+)
AI+,gCb-K1L713[[F@DVbMOYdVOYb&eF]8:/JgDcZ06Zd]5(+8b[,.B[e8@UE&HK
\L(XCDGgf\b6?3DWX3^[B]W8?KBJcQDaFEJI\(FJ<B:_/1Q]VUL[2/0L-7:/#:UW
9GYgCO\Q4A>adId+Z0N>&)^dO3^Q2C2K[C.\A,RD=+[<<_-CL<HXW]#QD/dX:JVf
1gD;Q8gBS30,g<[ST)@[ZQH-^6\=B-H968LYW#3Y+GI2=3:,<d0dE43SY@cR:MMD
&5,,#a\V>IfRGRE&(H;]<,@\R5(U/Y;,-J#VLQ8S^[dT5TgJYMUKI3.29XB.@KIg
NKDH0+L..QQLB]QLeX8f(S/3]:\0-KIO3db9=XKRRUZIP?1cFWIYW^)G+Sg9+?I9
Cf25.b8^+^M/g-2X#@d/ffYb12IBR0:;?G/R+,JQ+IBdS8cBHO()_UKN]/7UX.9Z
gI.R):6YZA4eZ)eN9]RS<EO<X(?>.K[)HT]?/;3INWH@(?g#.BF2L5b((f1(_EgN
W^+QWB3EfQ^CM_Tf#0A2>716N0a5WKE4LR(YO^;1/N<G=9YU>]>(Pd[ITfMCNQP7
:OANc_a-?gG+<9<M>L50Y=B22eZ5Y@2L)=5.RY@KH^Y:a>XHCg#9\cYH3022VPW\
bdf3>KW\<M#ZDA5>PVYG,bc6DdGcOEe_fXQP.>LL].cPOCPXf6CF4SY#ZCX-;L0.
eTR)6H_9SPN0)1;e&QN#4\K9#2>0,T+[Ra@).D,d8dJMa::LP1J)3.EJ<LGHC(,?
Hd.J/V16@bC)=C[]0<H4&^5S4?Ie5_V>0P9>RLR/Ec+AOBe>2b>Zfbd:Wdg^;(V9
NODCKX8/=9f]-Z>:FO+EK;V,9\49-2fVE)Wg,DfYM0.f@@LQEE+f)Y[,VN\9?3XM
;\XQQ1+8LFX,e@/4GNFfFDB/Y=XHNc3DBOa#Q?Sb?-=K_g;@R4P&<WWM:5._Q&@0
dQdM8c[46NYbe.=>6R7?bST;@>0N@;H(#TV_L&-=FB,?NVf4e&]#[A+ML2NL(KMG
6H/P:@4^[OX.dU7Zf]e]C#X=-Q,2^;Ie223g3510J\JP62DXMbfP6a/7F;4+^.>K
0+NLQf8A)EPT?D#?DH#B;Se0g-6&C>85)M&EQ+AY0_eL;5<H^./a2(D8g8N\,:UT
,H\:#.U:-]<[/B=B[L,>I)E+;(Z1;.(4L^-IJQb;#4(#AL<VW1,HV#?N8SC0>7@8
4TX\a>G1YX)bgbU\?.EWDBN,[3XbD,c<OKDRV7K__T7>@J9:J8OP,ZbSU(MaSg@J
3]LM>D<@NI@Q9-T,S0&E2AU<3+YE9Z<A_E<Rd?+)L1fA84#a3NB774>Z#HVPG0GO
O:-7KTA9M[AR6B9@P@BNTOFW_2R,Z.ZZ[AB+A=I]eKSJQK[K>]HMU\Kf::IW@;[)
BO3@BEJ]=-\UCZ>#3HDA8G)<+FE&^]a:;8deAD3RP99I(]]96=#N+]U+8P-9gSGO
BB:8bUKQ6+L+:3?,Yc?BaY;@)ME151;G9b@0=T7>G0-=HQ)d/FJRMK(+aF7D#Y2e
E.1gdSJ5C?RDT=MIP^H[U5U\+XfO]3739_P;a(7,bX39CEA8S5\,N006]d)>#0VL
]PaE\TZHe+8-)0_#M6:02JCfVLPD)R6&EBXWb>_9MaFc)O/&f.DfJ<N7>9a:PI;X
Z\4]I-OfXZ_;CI@+.AK]U9#8G6U/bfdRY^-VIIE0f:1#bV3VJ]cP^0OM@8R&K87,
0R?NH/V9R64b[UOGYPRV6Bd<_(5]d4Hc2NXLc6f0O7N3OP:>M6b[&CC9;d@[=NC#
,=?;&bPL1^WU3X&WIAIKWf0MgGYO#JbX6cdA1f)bW:P;?&CYg1YW.+3E08VS?4/P
D(TY6#9/\B+SUG:I5D\aZVR2>R[JILQ^?;<DO#U^RbPC?DZ]6[D+H)X,(U:7#Y2U
.>)La4CC.FdQJ8-]?<&5B7/+-L0-U?-;_R76@X]TYc^6/6/FF(UF\\/S(SA7O0bA
+\Tg@Pd=\]7@OH_BH:&W(b/8RN9?]bAa]X>CK;56X^I@7YB^9ER.LMAIEXT;4E7I
H\240a\Pb1@3b>A#\^REdQ[Uf>@A.+MB.[HKD?6_=f4(P&16)<W<Q:W/)Z<Z5@M:
?FEI#VAE7T<;=OZV>XW<)N-[EKN;N\GAIb-<9Xg0XXFWI8XEFJ3D-#/](IKDaQ?g
#K_L<#O+XAA>UD:4HZ5dF4ce>K<bXf,U;LCD8D^_N4)(U8SE596HJ9Za9L;5?A[b
D,6JaU5BOMcM]?2@fSJ0cBTF7:SB#[Sb>/b+f;S6fEEYBP]O,P0;0J?dad9U0XHJ
BUfC2@)8<@YgP&]+P3T6)WUL\8=@M,\A5cA#dH?4M4JdK78=#Y/?<:X2@bJb0RS/
,9-VY[bL_CJ[RI+-LOS)@63HdH^aXTKO:Jdca6:8HZ5/>6TfeX_+5IXGQR:PM)\.
;,UH(TS4a_58Q-1?M?S,/e=85FP3CP/5YYGaV[_=/VQg3N+DK@0_2(1QeQ@KRV31
-a82D;9@QY<R(Y[8X(;@)&c2(M8;W:&P_GcZ4+UN/)_ZfYEL71B6fQBb4QG>4B=@
J,\I2<cFdEd3Z]8GOJW].AS23eGY&3+<)CNF:+ZV8Cg#:7Ug^5O<S.R2[gHWeF/:
<FL7R\/TM+g2(UXAP;#XRT01QS]cIEF8]Z]cWLB94KU.2<b@WIa5-I/RKVd^;_?,
[?:S,^V1Lf3=T=PT&b4[\^.\_\U9E72>7B5.&R;JW0cTY1-PXQ(9?((AOCQQXQWa
1TLX2)c)?HGW86bOfeRN-LB3V<HYP\M#@H-^S#5Y4F;U.8<YNEb;.EAS3S2,T9@2
1RNP9C;fOZ+.>&A2.aQY:FVQ(ES/W<4[E46?]_5CY@@+-(],EYBfbVH+0/Fe?&.U
a-@R\4(U#Y]6.^F=:Z^;cQVT8G/^VX1+T<c6B;:e^bWU^dDTZgXC56P657+ISY@b
X[M6RM<MJMQW,Pb3(bVI@:f,Se9V<11=IZeF7X1-P.@414CdU]J^/A7]6,cX#eNH
KU58+TeOb-=,H74V9c>_,ZGFZB@>BU,V7,cc_1c/ZAN7Z.=EdO..U7bE/31(bWX\
7BYD/&ZBF-IC4V.],::Y38W7.EP;3]B\?Ke7d3CfMB\X1N(V#0C,_NDaR4?J[0af
^0IM=c\HTEd=NdX=[_4Vf2d\PV-0.C6/(359,DGL.Rf4I2#bK0gN&AE7EaVe:;Db
<3gS+.W_>L6KdA=5La;N=[e49?-d:K.UTSfQNN>L[R\FPO8,B5HFZT-VD=K[cU3;
7fcR#BF^LVOC:@Za>.I,c+EZ-=f7<I#B93S9Ac\5dGc(e?ULSN=gL?4C[N+Q:0DT
N\b:)Y>ACQP19[JTEKFXB<:0V)\Jce9L#b\c_20)c0+_NUHQAJZfe\57TJZ.3,O+
L/DV^<NATaBZ.SSY^^b#;Dd[UU@DKd8&bP4c;g2]F9X-+4Dd,;8cIEf4+54\W:-Y
IX_4^GD:bI,6ED\@Z(2\UHdNXJ36^gObRW]Le2]DdB&S,ZaTCb]6MX18UZ9#7-19
P[-41(F-0MKT7ZHd1^O8]eaV>),P\df^AB5Y6I<I^JPdf02[?:ca^X.M3UYN.DcX
]7aJPK+MSKFS>NOg[/_)(e=S2(JY\0+6A,?&JZU]N?\P_.TCTdY#KS(:^0RTPJBE
:O/4a5GD31WQ4]D,NLY8f1(>-.2gOD^Le>#Wc;/7V4^A)0?PLEKacB)]U3[CK=-5
YBS?:^Y->ZIUgK@R?[_4UeTN?0WJ9X:UFCHI,HEAB)76Q+DHd<\d4V)&?,ZZb8+<
+(abI;G><@1,PV:40B7W&9JQ<aS)@)gK).+CYD@FE/#1_JaVcW3BgHV0bM)f/E3F
MV=7cZ(TI9I\\TU1b6d^eRe_F-0eS3Wg8_)2H&/T+Q#B)g7N=GLe5MU.8?d#PZ95
^^.SK.U1dFA)&cGf8<_#aMa\](F[,GUWQ00A)A1A9U12M+8G+\.996<RO<X(c;N)
6;gY7X^fBba_eSbZ5e+5b1O]9SKa6798O0ZAK5DOUU1fQg\T]cAJ^G<:DY1+6Q1N
XCD+/(a1I/E#NNC#8BdWc70&8fJ[XRIgYEB[@d&0>/Tcd=(gEaS7RfS#S-<37.:A
,M_,REc;V8[:3<I>D[ROf>)?<2(9VJ@V>dKeOfX9FM;\d,(ZRJ,;5@7;ccMK48[D
MdXI<X=OX&SKW,Ve._41Fcbe(TMc1Z&M9[OUK]GLE:e4KcQ?\b0OI@KF<T3R5F/d
IJF52U<AS5C84>/M-UJXK;IN>RCK&Oab2]9L,\4e2bf(>F-=?MeLTA;V1S0:Q_g0
)0Qb;\NGT\?cI/76]Y9QcQH<XHWC,+a9@O8D27F0cc=+2A@>>L&Q))7C7[@O[+82
,1&.^_@QY-VQ1]UBa(aX;f;N7VJ/TcDP3AY]FW<f2UC9_9EP-JTMT.T2:fGc<@MU
>8U?#6KE]S6A9<#5_60TNN9eLV=(X9#)XTTV_JFOXMTd>-Qf]ce=gZ+f[8W>eK8]
Z:(^UY-0RG9Z)[-ZQW0@WDG>P29,B0:O85ea\DDL7Y7ML.]Pf&U32]]bM-MQGDV3
_Pd:b&5S?MP&^g9FfRA;&aM8HRAN08N5UJ38>\/:6([4^RR_0+@HW1==R5JNaXAR
_B^9:a:ETae\&^H>5^HV0]\W671/G#(PMBZEa1SORZ2;?5.0T=BWP]K?QeEP61<1
BWA>Nc&gQIf57UAW1#(JICHT]JNV&7.B7))IKQaB7G&;;IQ+8_Sdf4[J>N-(U<RT
IZD/3L)+9dFLM9S[](#,N+?.>?6WgB.;Z-c#OBZSE5\0;^XNL89:/P8+FQ[X42/A
:J412,EWV+aA71c3K1U+M=aeHGHX.1-LN;8=^T_+(Qb()>8ZX4##LT/070J,,:49
+a_0<F=c5P)Hg7&I(#KKK@NW,L_A.Q:e7=KMR7FYR8#=X-f.?e7YKTD^g4/W?G/E
]TQf[Od+;X74(S)d2DH9P;SZW\@,gA8V^ReNd,>E#g9LWL<beF#9XN0BF_BUIKRW
]c0b0(MeOIK]DNVWJW0&;CWK^gW_[]+D#>P&<&ZI;Y;E4C>aJ]>&FLgN-3PP\HF&
fA.;YIc3QQP7#Vf.6cb.?>G=9N4Q9O5Ug^1e><6e_U45+.,L_S_)@Q0<8E^dQLG5
L(DHZ3SY-gJ5T</)S-9g_:c^W?f-@A^b88@SN-KIL>MNKN9dYI)F56D8SS&S.0,K
EeK=REP5dF]Ca_3>A8TIEMgI\d1MU8[0]9Ia&[_;#K9F2XP0_99bXV(CPS:3HPE:
E.GX9IV&L-+fB_74\B#K)XUb&_WQ<3C?Q82[T)5GMOdWNg=fE0)P&JRcE3RFJS,f
V])M.EROGT+I8E6&62Y2XKRT5I)HE=:F\A8IME0L;>C[QN>e4P&JK+Y:XN3GE8a6
M),[K<a;U?F-(A/[OgD)7+YaFO_Be@<S.86&J35OOQE[DD/:UVX68]TK0#_L2KP2
.c,]<1&)a^].5_B5Q97eGH\dFK8a7@9TeR=O@@CLbQJ(V#(DUQN.1KM3U-BCgg<\
7I<EOV(ADT:]JZ/XFM_G,O+KG<\QAe0UW[EO9W0<DV:BJbKacHC\50+KV>:g-U@+
g()EKf:\I,OOdK_b^M=Q.TGTVJS<)[4+9W62<D:XN4\cX?=4^CeK7E2HQe@GFGT[
&@cRFMB.YD^&]WPV+Q.6:CaPLWYG]J[=,9/(g;f6X:XL#SM1O1)c8BCef154JeYA
A;9R@&@>#XG19LCg4V=^3G\c:&FBeE]?;:-72ADd<fI[3D]OK(Z--R8d=3M_W#);
)PLE?76UDT0@2LYN-LT/)M-;0E.#KdW]JeR<-S0\gbTV)(DN(0=\)#5>\0,^5JXc
9.@O90)gWFgODPY-I@d6OO(B(bHBFaS-EPJd:OT7H4,IM_A?<JZ2=8<</03Xd>(8
Y^-a]=8F.,__&K\IK_R0U&6N8L9V3O:g?;8FW@Ua^bf6^AOEbMP@^T^4B.6)=@8A
Y>LSL3J)bbY?0HfGT@JHI8DUXI.V^9eW2T;JI7cLa3\<TAd3@>S.:4NOEUHC(E+A
4U70,#e2HbX4@9E=V)Le+@=@8+C.F,V/5M4)NEL;^30f&0-+@&[^AHGRY2KO7MP2
90(EDaVI-Ke1PKU.Ga[+S2df3PR7EKRdPBe[M6:I_JU-E,EGVWFNB/PS:Be6AY1]
_5A3^P:2V1?TEOd>(J+gE^IFEUECa9+>dGRF-)Q]@f7L]X+[b-8ZB1f?;^R&SXRD
fRI[aE_WIMKAR6a0#@SD86_@S]8;e#.XC=V[;>3@2dSPe-=+e&6<cAV3JPg6PcWI
)1<55A0MI#L>N91Y::?\O8X\N0D/b^Ma_gZH7fGeEXc_B:[4W-6@@&A#HT>.N,>:
B_]PO;/6=Qb]6G,2C=3(=E>GUb[JcRFBTIJ(N6&ZIWZH(5[gC,::ecbA_CdUcb&E
T8AP]e8S_9Kg3A/9Z8fb@:?W//T>:5d7(6C2fbC/ZPOfC)TP(@/\K2IHf@D[JNXe
]dCXY]<ZUDcADaI:Df-IcUX#SWM,(:LJKda3Z&);L6IT5LY]M1E^VZ1]Y@F;E7Z_
B+=FQeNJ6eNTTXLO_4&(4@RLX3HeN6HX^P7=Y<;?CQ-MT0g)Y>_EF.OILa<36)72
[UH7KB@Y35<]bf:FYfYT>=-/LfAV)QM-5fdY9Yg/<aO/@#O+78G0TGY_ODATE_1J
<_;e30EQQC<0Y;cI:\@D]eE6?bbg#eC:F;eQ@SbI\QS_1.c^[Y9-.V8[B_H]a4TO
],fE;]V/><JF9.CEUN5JcbOd&L)cC:cF[ZGcCO]c]cDDT\b.W0JC[Ub#<QJbPIAW
f8Md_2.g?62MeS\FXHgIUA5:Pf1GdNK4PTVNc(ITEQ-a<b0?fAf#RX,0<MI7S\Ld
^C9OS7;^U75:O>R:;/CXOKFTA+5&(O7V<[&UC#<&9O^Q9:N[UHA@&&+G0acJRN8[
&M_PNAK:M96&((#Cb1=dd[7Dc,W@N4]TZ9TVAWc40>8/_)0Q0:#A7P-,H>54gWJYU$
`endprotected
endmodule

