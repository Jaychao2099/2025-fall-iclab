//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2025 Fall
//   Lab05 Exercise		: H.264 Prediction and Transform Engine (HLPTE)
//   Author     		: Bang-Yuan Xiao (xuan95732@gmail.com)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : V1.1 (Release Date: 2025-10)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################


`define CYCLE_TIME  14.2
`define PATNUM      20
`define SEED        86

module PATTERN(
    // output signals
    clk,
    rst_n,
    in_valid_data,
    in_valid_param,
    
    data,
	index,
	mode,
    QP,
	
    // input signals
    out_valid,
    out_value
);


`protected
U[1.aOUa^^BN<(0GO,YQbNEdKX,Z6XQI7/CY(V3[B+YfZ_@C8+)U2)R1C\Ua:F<>
gQM=#a23dLLA2fg9<LBLd.R?#8\<gbd(?8]Had83/@TfW@7.C_S:OHD=7\5Ac-(G
3461)d4T7]&F-:>/R.D(V#H(KY4ABGF[WcMD5VE&e(6d,,J8K80#AN1G(g]6a9e(
CS1fG=7J)32cACNNSWP^-UdL.eY]C_OJ@^NfP3fKMR\dA$
`endprotected
output reg         clk;
output reg         rst_n;
output reg         in_valid_data;
output reg         in_valid_param;

output reg [7:0]   data;
output reg [3:0]   index;
output reg         mode;
output reg [4:0]   QP;


`protected
A0D^WH>J5Q:FQENQ=7PKALa]GbQFPcg1@,[]Qe90b;[&[,V_6QJ@4)eC6]4+2?Xc
ZPCK]/&e+.T5-/]VS6-&aKa]2$
`endprotected
input              out_valid;
input signed [31:0]  out_value;


`protected
4+/17?)Qb/S?TNNPAVa:X#N/A]<O?RHL&,<XI.SI_)U-fZ1N78?,+)^eP1K_ACDD
JLZ]MC3;N0?1U-?S3^@,^8>HAS,.EAXWSO\;51(SfDdIQ.L-NeXbB=VW-M7=J_Zd
3WJ91+^KL5J,PQ0B+<B-XJQf9c/8Wg4eX3+(OaN@<-LL&<]ML\<cA?\8g=0[Nc0e
Q\WFNM5K6:P29/f(MI.BGOeG9KRadf9-M(PKA:Pg@SXL)7?e>##D[f&G-Paf6CXO
\af#Je2AE]W_:_F1^aPN1]O1A9b2c9b[d/X4(\1N:(cUfQUO]8P/d521)N&9&WVd
[8ES\(_:1eI7KXXB/V\-gUJDJ@,Gd?3B+F)7\&..I_g-VHC#FX5F@Z)<PSTE6)M#
Y_(a:VE.X]0;_?:<:V)0dJGJ&>&VL80(]>WDQNG[XS.7JV)2E:(36GQ8b0,&9EY]
dSBDXC]^AF&\0XPWe5=J:5C>3HV_;-[T\QP;8)/U8P?(]&IH?+>766SE9H9>e:E/
,;Bfe1aWF-6=g#G^VaI.,SW]F.N[Y@5@GIV_^TOKJb1J7&@N,JJS6LJ?1=?A,<4c
^bZKcN9=-?)-]@&0?Af.b:3.:CfgT44;4PPGO2U1CR3MI&9/<d(bC1S[YVWED-U6
B#dRU<YNd.YMfAc^CRW29\R<[X=E-cA)gK0PN?@5F&#:ggFY06?,@[<HLf[OgBdI
>BJf&R6NAQ11;L-,T6\_G)gf6M-TfL[aQ+R6EIVZb]:abB-KO<8Gg<7e-XZJWM.,
5G;7=NdSW77)^2R1WgRZV^d)KB>V,+326GTWS;Af(PE5L)V>g(/K0N+>/g(R7#?@
Y;aMcgZX/gI\EQd:+KCRE&]Q7,]Cc4^G=CT=H6Tg,RS)bY^H?6?U#PZ.JK\,/[BY
N<aDU<H8&71><KJQaI2@QV5H)a0B=&Z=8BKL3\b(G(4a&UgR+39.eO?TO_5A-M6Q
L:c7=e4961S2#BC+G<RZ8Ed-O-Z;B\,=g/]+I^]MH9gVUM,T-]0&H@T]-A)^WY3L
_[>Cf&11fT@RXBg^<LQ7A4)Z:\_AI58\T;SI):R,V[+M>S+GTAG]JcVL.2C#4:I7
V\JcE+S\b61]CCH_=WLU;T@d;b#(afW?_>6EP^;<dZ(-&K&Q0/<,W(DC5)MD/;H_
YSYUgLZETB9<//FfVJ+];VZ5:@ZSR\T82JfP^0G:Sd7_(A:TUC\^0TT?,8OTX/HN
9.U,<B>##H])K^d5UV\ASS<4=8TM_96>_9GDb\Z>>G^JD#USUOZZHdA=JQXQ@c3?
NgaLZ=K]@W:GQT7PD9Ac];>(Q)^cC.[2.EA/J32b]_:<eDD@L=WM64V+bA<HYEU@
]=@aD9<27@BOXaB?K:NT\_;&V_=IFYI15U6M4QSDJZ,>0T4g7c)<#5:A)HYMaJ=,
U7G@Wf)dB7eM4HA;Kb#g.VH0-)<dG+9H=QOe>>I65\TG0[6@T7c;D.8c:1\TJXg5
8P0\^1d24CbC&O)_Yc>Ga9NWV39^MR3)g^LG_bG<Wg1eG=FFPC5GOXMX1WcK?IID
^gaR&A7_S@V>^agV2Ac1&ReHG;I,>HK@Oe7#H2(0>4#9?DKCV[B@@6Q^&>PU-U7^
V>/,\>?<OL>[f^ed@;B<XC3L)+Q8A4@<<(0-W?/<J07gTTN=@,89SJeUP(d-)fb3
b]d1)Qb9C9f4f0A>(abVGJbT;ZBg.f]+?b5YcH(6fL\7HAb+Z#CP[&GPJMX<-MLC
1VEU#\M7TVCbU>H#[;EZ9194J8_f<^HBbe25&\2Y8R2W?Jg&+_U@NRK<53..UN0e
B;6[Pf;1gGa(;8PDeI_+Q,079;4=L.#2/Z>,LcaVUS<INe?b<7[[)@06O3_C>BSN
[M,W5cNP:58K&&N5\6HaZS3[#bMP+FYO2(_DTZ],N(<PJKEN95.SCTN_,7C)XF1J
G5?ZE72P0NNcH\I^T9H#T+S/W&F:bBU8_Y6>=\g^UT.PPRF]=J;V_R]fe9ebQ8^A
J5<=TS_O)JI@8)S##?J:(\Cb+9_=QHHda>+9MMMKC=W5JQ73.XeE&_O1eM+)SL_&
?fO1<\E^-,WBd4K]]&1D)2KX+=U.RJP+b\N2EW&21@:90(I0-XCT]52,G5NR/\-R
&A]8VT/Uc1NAZG0ef,&Y?0KTQT+eB;:F0[_BCX&QD]df9>\AObW1g.SZKJ4(2N\N
Z?:A^ROUPEAN^A/1BM?>4c^111WD6SdM+S,7H,+C1YK.5<?=#aM9)>YD[9Z-F<1,
.=WD^EO7#7(9^\dVN0fSAH3N^dcYM@(3b/]3K<IXO1\VBAgMT92D)b]KK(^W7.[]
AegYaCdL7:,)-U<NBQbVC)V:BX>N,^/6//3AaJY)CcDC]07g0_AS74dC64U.cQf]
D2QB@1QVBXHAN[f8VR\F0]YQ?O4_9&]MMI,V23eXO/bTAPS=SK>O1LLJB@PCaCdI
5]GCS[a3fc_WB^J1AG]O-=dW/@Ne#dRYeUK1#DI#;&,<-6_Y,D<-0R(?^dOG7#Ha
8Wf05D#]cZ)/SNI<;:1[I5fa=+#J_5)I)A+H0JBb]X@?GHaH_GBaZ+B=W)/Q&V[1
63G=I=DYK7^,)g[(^;6?V/P+_[H)^CTV-/^[I?CJLN<F+#F9EU40\\K@c\UX[0\6
@eeW#dfUDT,=P1R/SeLN0NBdMdU\(28XMbKGeC2]G\O[S-BV2A0GB;V>cODMEQD_
O)@PZ#9RbQH3.G4QV-39JC66>V_CM1gG;)99>MK2#P[5b+)B-K?:5,a0/3J,1eED
c0Da&-KG5dXJ:cB:<Q./(ePGcV-5.N;efL7aG<UIVL6);[XYU65;KDOUWV[04FK=
L2,WJgE;.]d[_6-P1e0YFAU.GY\8b;b-<&=a@6[^BL>^#6]a@6K0.[(bP6<<R&_7
abULOHf+\+Te3Q>b+#S0OH5MD15>A8C(]YVSRF7G+6>>^B89f#(VTVB+,6Ff_-,#
5F90a)bF8)f_^I4PU]:#0AMQ#2=<a)V9))E7/MJZTP/L6D/f,N]X.=J,/2Ve)DQ^
WXQbOJ4:;2+/NYA,^Lc4MWI]#H_&f,,EI8K#8&42S+Z-RYaQEV<>=R+E#J3H;WDb
D+BT/e\,\O/Ebef_V.THVY3X6:&7A?dG(g?457#(\L0L>BO5;:6E\MNQP(8CBM,[
VNc1KO=9cg^H8^G-c7>eb^#C>#Y<^Rb9?dbPcM+\=J&E//.O2-_6PT](R6aG(S7P
E6O[SH8R=7WY3]<\5HME9DYK8,)7J.[5aG&;LGXcb5>\EZ-W2]B6(N7:5(<35_gH
J6+7\RH0LGEJQCG,]@]4]aW0J.8D;DSB&6G?,34\6XE<eJ4ZWN&?cW#e)N+>N1B-
3:@)0gf7,\PLK=YNA@I+S02)]M+>38NX973.28_5#S2O3R0,I_65S^B,X=K&&(Q8
/:GWWYP0^06XVfbXVS:ANY\,;#HV-6W>&83S4XHA[X@YAOL[X^((5Z8D+VMT?@4:
I(YF(8?L>KN\X+]N;(M+L73OHeR]?^).=;@F99(QaV&7]gG#@Bc8J(0@XOG2MF=J
e.^G]RM=RV5D0.I82FHHR0WB^E(WK2Nf8CL[[GJ3T7&7D6N/e\]cS?)(O?<#AG7Q
dA?<YTRYD(JYU&O-:\4K8:gASOTKX[K3]8_Ug88)ZWHXdB>DF+C/dD?aM^Y>6;RG
UU]T&N.IX28d;RLS]S)]Oe4X5^W:]>=8BcWHaC3T.+2B?d)cgCF=3RO4OSHK(\T4
5Oa&fB.eD.d+@M/+H=.5A[\JbRYZPd.4Gge.N58[ERH7.#M.I>2S-HDeLb^U#8ZB
SALeg-Jc-L_(G=825HTf@#^gF-+6.=##(dB2d_aacR79gVH)N.,fg3;(KS_]>H8H
HKIHP)ULf;f8.;a5K2[,\L/Lec.L1a5>02NT\5F77PbON?DB67&>?J^,Y)M]+?IO
b_S8P^6VFTYNKE==B?I2e4M:<fd]QP>WNY_FMOe=HICS3O8<[Q?K@^N@FF6>B6&P
6S195VO:)6&Q\P792,#WLEYdA_KgEGCb8Q_-K)BgME+R<aY9?>UN6XJ:</RW5>/B
_c6#23-WM5)-AHJ/17?MGFeG6_R,/<#;b(ZBd/@.-98/UC6710Z;#;L>VQfdAZeM
9+.2\8&84XH1Q5?G\>eUC_\N.7I7=9OSJ@UaU\9fO\+QMc040\5KG<7DZ/0BA-3d
g\F\8c8A<]6KT-R&B^(:#Y]<,QQ^[(JEeW0fAF;RGPc]-=<B#f]W((CHQ-Y4e=a_
M@[DX<,XSLZ?2)d]a64/H&5PK83&]9=?C0]7YAB\A(52(-H.EXZ]V-GVP,W57c?#
e&6VS&/65#;MRUaa,^&JWF4M_)(UOQJ8O)H_fFd:TZ/Q+P^V1b_5/D+C<.;6AR:,
a0=REM?YQ2]26B^6aA75Z@:c:QeQ^EMWaH:]IV.A\4,5^M7VTB#2JCP)_X+P6XdL
9#Q-^4=G[2UMK&<../Bc?QP=Fd)X[7)B=/:.X<F>.??K^.^6RR72X-0bc-V/QGR.
ZI1O?KQ39U71-aaI>Sc/NKP.AZI^J@-(S_F^7_=#LE=geTJOZDa/eFb[?3Z&N\Ed
STC-;,bF3>/a##H9K59_d9eH+d)2OCPOU8]6PZ_9Ug3gIJJ3GR3\dA<(YFWBO/#8
)WAcee<?IR.=9(4S&Q8]e@-K)dF(./8_Ne9J,a;cK3J]U_fX>HU:@2W,8;1;ab5g
FSd4?(UP3T&31gBg-Z^NUZ)8Y4\O)f1NBaKZM0T4f&#GNd#C\5#-7;43G5/H0&e@
O5_MLE6BV(9gJ&?T<68@d@,IDM7^ES\[&,XDYPa_f4YSEWWA#dfcP:AB/fAaH@F]
WH3TMc/WN,?KFY/MMe[WD#/0BM59[<CSUEZW4@GaT9Kc&+B1P\;OXC(FBeN_cc@L
WRe_dQD=O@/dO,746eRK)YV7>4XC7#d)b-2g=9A0I>HN86dY5:Q/0^a-U;F8]@Z5
f5ODFf6V;NRQJS9Z8A>^G4>E=X#/M9P<f_G,9S[CDFEW7LRTE#G/B.>4dUb+[,c>
b8U/fg7bOgP,W&CHO(Q7bY/]B6RVR6Obf+CEW8B1<88H.SGE#a#(2EJ>#M.\^aW?
.&U^cA]:Je-UZG-b5bLB+^c4K<AQ>BK?INf_-f8A8JS8P.1UG/FY]>:+?ag0[@Rc
F./DNJNTB3@1X/45/>FgSM12dX_;O0b0EV)a1&Wg0S[c,5_cKI@OU?^]6BZ^c4&H
/6P7Z.:Ia7+S9g/4KcAaA[23S5Q/UB3U?XR&:K>1<<6]MeKNVA\f(:RD/6IDDU/g
TU;@YM.CS<Mc8B&H7,G2T+DOH+c]I?=M<:cQGD<]ZOVYEIfO/9<LVEB_DVbbBHT#
A091NK3bR>V3J)\5L3OW:&XFf^#L^;b@O,5(0KD_:(EVV@OTOL:?>e5T.2@/M4&9
+RK7CeJ3<_VT:0)NE8+=N?eSHfZL7&MB#[Z\N_,&<Y-(TGWEb:[F#<?8(]N.B)TH
LbZRT75aEJdPO1)e:\;0-2@PLF(8C1=N.)^-d@[X/?#Q[C>Y4_Z>M5N8^KG;6S5O
5M:A[SQ@29]fCLW1AYL4^]E/b\a_fRA<cEN8HUW\cG])5YG&3HT(78J\JYEb1:9O
](I<TGCa:;M;EUdO\,@R,P+&S2LDB.[gV7#1IQ=Q7?c(H3W;NTKYddaYZNQ@60KE
S\e0;Rf[+2@?/\H(,7CbbfGb(6YT9FCg^IH,UC.=;YcY7B<KXH-EIQ7_MSBf-[fN
-1<P?)RKbQ/_bg^fH?C-8c:HTZX\>>86=TIMbSDR/F<b<RGD9EIB>^_2Cg-LX+G4
H4J>7^B(VNW2&D[\Z2N+adFC9,[7_N-<-M7Y]KMCXdcZUYacT2;2I@Je4[bODGOF
2[X,L;a\-UZ2H>POg1CNAAZE,R7I8KZN2RGb=FMf0a,a?bM2-K1ZP0BID7LVI:=c
5E=HgVC>aY?;0fbIX.S:K,+.7:7;VQBA3]Hb\[]F?J@L[U(90[cECD=R)cL7T#cL
\G,gb:(L,.:ORW39&aNCN7S+J5-f86G8@4GU_,7R3+[,Tc?\WW]5/:NNZN1][BOE
7#J@?0Ua(^D2CfNWe)5G-0Z.)^51)RHTNbH_ATWD=\+EeU;bS]2(MRQP\eDXZHLR
&.:-.82;?RPF.)D[^bIP,,.6O[7Q]TA#>T.QLZA&Te?T9LdB@...HBe83DAcdZHL
F&,R[A,?D+^-8bQ6_/g;Y@NO)2DN7R[6#eIR\9JZ_d_:\e=WIOE(EO(P(WBaOGXY
Lb395-73c[aLTb&TIJb6;cRBY3DQ&K>Q2#fS^?d@,U55CRaVe<C7eMW6DMI(>6.U
Z\(YL5BY/6IfB,DgV94+1]<RCMALT9?)\=B2R#;@B#+#Z0]cfG[SX8c6)KJ+?Y(E
22:1J27S:g.Sb#g3b8?DV4MRJ+15aEFE78e.g&C((_QP-IgD3FJ5PZ5K+,MO_9WZ
Ja/;Y)&3ATAKZF.47].I1V:A9.W:D#9?6-d:K>_K,NM?-^FQ]1D>G#O8:]-C8.1P
=0R(0b5^4DVQCC2Q6/:;:7LFf@5dQS1@Y>bG#M#ag5TPC8Tg_Z_HN0QNd^=XaJQ]
+f\2+M5+d_G3bb]g?VMT1f?>+56fL=65\\QN3d?+C:@2X,9G^(5<:dJOW7O/C3?C
@&AEA(f@O?_M)/)+&PTZQ;Q/8=[L6#;?UR0X<2RT[a?Gf]RKD6UEPf>If))X\DOP
)Ke[DL1fP=G5U8AUZ&H]SbYI><]#cKg8E]URd&7LWd7Kd6-b,S1SAHHg^febXP/C
56&LR1a[GL@##KHJg)?U-^>.@(>a8<^^RZ;S42R]\^Q<O.=EBS?Og#=UAN@#UbU=
YLIE_HJ&KO)<=+CC:;<2aM8CD:DNB&I9Y>N0TA8RZO6S69JJ?NSeCR7+/<E4B)4=
\>HO(KeOW9g07HT6P#:<3.IS(HHP6H[.H>E8,0YV\Reg@F++PTYCHCa#-T-<<dDQ
gS7@?=6CBXE34OLW-V:B:VBf8=)?P=GPG5Ed(YA=g/62::NN[C.dWC:eR&UB;5#W
=#f:eB8B<+D_MTTF4B;M-d?#I9>9GX4/.YH^VVDO[dU^6./11EXXHF&D,L,(3U_(
DBdY:I9^c[#W<D?c2Dd3#a7#Lf_Bb;^,UaI>4&+g?P.[#O1TeAD]W#)F5SbC>SY;
F=@K=9YKFABV+X?(B(I3Z/UV]=M[TB>YH9T8AdMZY(ZN5KZ+a8VJV]LCg+4Q^QH3
<fYJJFK&C?:2E/,-0P3Y5[HERJUSX(Z-#(5cT8TAPL?KK,fR2\[XJ4GWD@7C;N(O
Gfe8HRIRHH:IC>)2?c6faTHbIO7<f6CXgAE/V]RIbI65+M-<Dd;D4-_#SHNI3X1.
g-^Y<g#(5ZH1D@d>#14S6O[b#]6^+SREIL9#</S>0P/gE1acBL&V]e>9X\_\OJaU
QI9NL=f+LMOGQ_&aae+HU7)\bYF(=LCL./-7WLO3,BTd?c[>7353L<JgX=U>Oe.N
e1E,RgJM),][6Y;Qdg>R?\6V2Y6[?3GZSFe58;YT=71=O_5DAO9K7EKF1K=T_L,Q
d7&Z#)SbJa&C_=XB;I&<aP2R)E>]Z5L@[:);6:&ZU1HJga\O^(LX+72Z/Q9:&a#X
40BbN+:LgDKa.N6TL^&PFF[=\F0V<V:U8MCN6T@3de)c34MD>_#_RQd-c7R8Q;C\
aC_V=5TC68AfG8)1T>^dU;BAMTC&Fc-5aML/<<],Kaf.]\4E&[GcXbWaN8EW?/4a
,DES:d652_4c@ADKDZ^Nd-LKOY@G0^5A.A^e(NTD8.;LBR3?0(X\>?g,c,_Z4(#^
=Q>W5IWM2[gTf[2G5I<VB][\0YDe<K96>BS2Oa;=H^@A3^0RJMaL>6ZL#_Q6(::?
>(GS8Ie2S62I@;8@KZ(PW_,5(@?=I?V+U#Y=VVD+ANO<-^9aOE>e@CW7dV>TMCYc
7H5egZU1C3eC?:E-N\6MH(MDGM8^6&]_Z//8M=<O?+#]NT7d9F46,8Uf]e/L._7[
\>@>\8]I=:3<S>VCP5;.Z2VNY:S6d9=:+Ke&SZfG[5dAL9.J1=><NMf0FZ]+I2P5
c3Y=MFU02PQ7Y]-G=2E^XPT=@J24VM(T1.>NYBMVRZWS+1QH;_PZe+NX=MZ5S8Qb
Y9^0JGT.GB6#H5IB]?Mdg-(XL)2/N#_X;O6IS>7W8dK>9=7Q0XA@?#&:MbV-1If,
S<8L5aQMc&37+GB;C&Qf;0KMY7.T60C^f;87Q;_XYI1\GPCDZ6SPfgFU5G_edg<A
GB5bT2H>/,FY77JTFT6WE:Nf9D[_:3V#F-=&WL^D:VV3Oe+UI9b9F6NBLX78c]9f
4.B>SBg88MN.39)4H&7Y+cT6Vfda6IY)gNWDJS;b]Q9W(HCeSd+HIg9C)EC^ATGO
[#=ECE00NfaD^HXS+9NBGeg0[=A>)JB&F-_#P2M,5&5[P5/6aHT1L94CM&WPD;/9
TRc3_54D]C86<eEaG:.[.&6?&FTa(CK,NDCAa[/3#=9:-#Q3BRM4E@1;.RU/?<<.
DUA1[N@OU?,49I=9=2ZP1=fA)+R;=@RO-IB64.bYe.TN_1[67)C==:[MAfB/:gIK
TGC;#fQ+MTSO)7cC>-#7CYTL8I9<)H3:a.Q0RN-3TUE;GeFA+GG2[=HPARJHMRX6
06dI+P/a3>cW)2QJ7N#HK7@W_6ASaP@0RO^)@OWeRT&9L9TXQVR+J@V=B@6;N3Xe
TW)L/&V;Z7fbZ\\J4CYG:@6ZW5LP]gcJ2\0.\\Q,&8K,\GB1e;ST9gF]>(B>WA(a
#;2@R2F2RM]I1#,E(@_/5K\WN,eA^NS),CHG-W;E<A5dR^@N[aS^d-7W,Q46:f?W
5A&cZfO3(@a);WZfSG43Z/N935;e3J^R7](7GU(FY<e_C>VQ_6cMT.R(+0D7Z^.X
&5=8>(Cc1V9#2TD7ST##:#;Fb/Cc(c3D3XI7/2Y9F)7ZR9WKWJ3J4N^BHEQW<Wf#
)O+[6R\#O?/B;.X-1UGa(I15^3^N)/GB.\T.dJ#&B6L5Xa.^^CHaPZUO\X)d.>1]
BAMd?ZUdIffCb@AJ#RQ[79)HOB8@gQDQU-;d7@^05=9aHeJae7\CJ-^LRP=O=/]3
X48(RG\V25bK=NXS=\#DN3E6OWf,S89XLLKT6P_S6KL=FG?eTVFgLY5>&)?J2T#a
MHZ&&2W?4<QZODXNR?PU6e(VJ53K@.#_PP9A(V8AcZ>LO3Y\bZ7KQ]YcXD+Q^cfV
ZAf:^T]g^KX8BF_BE=NG=\4eIV91g<\>C6>a.DGe(FaNPa(&MT@^#Y,;GUe:&U-6
<:EOX3BH[SAV:5+H[a[50>NJH;6P156T>NT9FYd]ENLKDT>YXNV&]__>XJXbGJ)Z
WHM;=-\2(YL;GXJ1P&aU3A,Y2;b@L4PN;F7&9I\T14g_H(6+E]J(ZQYI.L;@66<Q
HF]#C=OdM\LX7E[8/S&R9#B5Q+E]d/:O:a/:/MJ;G=69(-c-W[T353CE<1bQ;4bf
CP#e?6cVQcGRW;-)AA^CMc8KaH5FL?@NB)QO=0SHYd8Q<Y36fKS][UDSM,+Y&@X;
GFRedg_FFHRd5SZK@c-.(R>7S/@/]D6QY>]aHY+6:>AL:WC(:J4N0GFVTK6;GCAX
SCea7(I.7<[I=3?Af5GN<aaMT0#WF+#X]eS+(EBNcUGG9/<8;;[PWPggT<@;TDJN
#E(E)LJWXG/)5YW-\79:UA,_75_A5?S]@3::aZP05g@3I50\d?AQ)O>J63LDU+9&
EB[+aOfLP(K\L\<bI6:WMS,5T#P-SBWJUQTSS1(ST#O<CA:I1F,d))VYPHQOI>:2
E+VY:1^>@J::I/MK[eN(MJ]\@DP2gESdG/5#,U]D8bg0?gK;,N\K,T>OP?].X:VB
K.W++a;+f><CQ1UGfDR1IJIRBRbVc6CX2ET7\0/S?Q)aP6TL=X-&>B;7C#FSL7(X
BL;dBW>V,<RE.5<N?K]52R2TK0#ZA4N:\bE3YYV0>Y11OK_,L19a(7F6[6TX(X.>
=]5O,I&N&37?Q)_]46>IU<C?VCZ,c59)<XXMMWXH(#GZM\?,KL^QM;H?>L>#[bB4
-b8+]\F29bI)>ae&F3F@A3Mf5)We96Ac)+L3Q7D1gS>,N,;aWR.Q(_IHFTMXSFLN
9BG01W/Z_)eCgTTROMc]K&bIDVL^N&fVJUD&c=^Qe=A7c0_=:1EQ2a?LK8>>2/-O
BK.18f\^#@#P2C\]@G0NaOeV,ZU//d^X=R@e->LBXYd,JI1<<MA>S;5]-EGFV5-A
\+bW3<g.7X9@7\((>(DHFgB6HAD409CFgY88g#=9/.26:2MF&>6^DY/MW@@XJ2M7
74\_=3bcYX<FE:9/K[T2db>0cC11R8<[\f,J@VXLg.:WZ(I[;37[]([D#;)O,[Uf
)c5/JHH..E9b#dPBS]WO.C]@-;#V_Tc@L0(cdN?,E&\JY064HN3NS2_FB+RTNT]M
?36?FHJT3MbRMK.XHTE>I90gU;@V)<5/aDIKe[+CKNS4-9gNZbNBSf;gZ:MO9c\)
4I0T&9,aJ(e>[K?Q7-F7MP82<#PRdX8<^2H[4:57=9B=/JFgCVM\/4_,#/7Fb0Y]
AeI<5YRY;0ISdL)N>e<KTUV+):Yd1YKdc;]Wf=41X-Yd\WBE&^6A0G_S=XcHP,A_
)F6O2L#RGe3WG[d+0]UZ_F/1BKVVc5(f]fb=)PVPO56(31,N5SH#+\1GL#2aU>@T
B1P_]-H+a6W=]&e>+R#F1bS98]W6bH:<+CD5IR--K(>E8X/DIA.Z_@KY<&-K^aC)
ea(cc]_(/044A57OUR1acAPgI/;KF9P9a^2J[\gXT;eS&SMdP;c69)O4=dE,EDN<
9(&H\)fT3RF^#M(=>?P#P?H+C9R7#7E=@SHg8a7.d1aV#[?#Ad?L/GP5Z:KT,6A,
BfPAO7/P5RdFgX#EF[/(5^,P^^T2Kc_g^JWd@6WBT6V&Y?3\5,+^:V0VUd>P+:W)
,dU/D;K9f\PcI-Z3B1<+W(C7Kga47466]UgTI.cRJO67Bb(=E/O?C=1BT5S@+U(@
?8,6@=<,JQN^BOd2@>LB^eb3C:e3V[Da=c[_0K_]b2GYaQ,gJXMTP?I4=2==)R/D
:=IBU0UA0R>F::DbK&CTKK@-&AdLN-C:#0,E<[75I=b?XD^G,=DF37cU3RA4P_RM
@WcYW:Q4?#;:,5+4CS]SY<G(T7ggQ&Z3TIb<Y#dJb7T10>aWfNgA#)Z,TXJ3>[G.
IO6bT6FLDUg&PBAAe>=NVTI+]MICV5f9eg-;>G]d7/]_F3:eKY:Xe(X2\0ZMf)^6
Mf/9#NH8?YY<a0?1Nb+-<IF)E6;8.;TP+5WLU^[1H#-EYeaPR<_^>,I^@f^YU==-
:Y<N;[W:Zg:,cLO:Aa97UNSS&gU@2WLMY.1X)56OLRCZ8-EPK?_M6-5/MF\UYbG1
G9(R4T8+_1#gGLJ+W8QceBcR2H;U>QQ[OMX@+AZ_L-ZEJcQ?Sf2NW)-^OJ[1.7N+
A>5UHV/)XN^5/?)7VB,PF,\_da&FAJ<[L:33^Te),MGR5@DWS4>/c/=aK5A?N#gB
=IEVGa6KYG7Z&fQC?I&2J_PI(2aQ?Ed7WF>8;+>DN8:C/<D9\GFD\83E,MH#W9M<
,00AT6JTUbVHS1N&JVZKP7b[Xb]]0</cQHa^f+Y>Q,_5b5Ggd-(KOQUCFOgT&8(;
(+^6QPB@UH+HOV9N/#Z^gIVFD>BgaUZ,5-/OEe9#;V^E[Z_.aa=:6bX=^7RUS0SP
3/SEMS0F3T4+B_7[_3UbfZW75=\b9P^I_?+&65MRM7W/B:(<DB:EN[V8f/gW=3BE
d@N4X@(XX2[b_CPZM=8He]:dCCY56&K:LIST6&S0e+K?3VC3DW9IT9A(g?J;G:NI
[H:#+)^C/+a(L9.=C14\@[((W4YK3J47JN>M0BFIC;Z]RBOa[ULZ=I_O9aR3c+NE
U#V\#bWQ/e6g/.^d7-_SJW0R:P00\&>8eA_EKf2O:\AG1c7P(d[A56W.ZP&#WE_Z
HPK&gf:T+NG4STFDC8B@I/IHJZS0^I6SGK1\17=MRd5G19T+1#P/TX5NNXbIFW@^
bGETf2&_8B?T:2a9;>gB6@JP2ZUU0gZ,aCN,/^(]#CMfGa90D,JfC#GD0V<X4JVg
.]K/bN=KD#ZMKbF,e,E4bJ1AWF@LI&N7:I<T,#(3+=53)ZA8\M(_]_=<H#[V#YR&
=\aOCdS?L9OOMdUROZJ2Lbb0c/+b<(H1VO3>Y&^7Yb)CXMGE?TD5IOFPIVFe_R[L
H[+EGDF>6X-F5GK_fRFgG]1>cbE]FB-M7(RF4?(?#gG-:O[J9NL0Sc\Ec+YN8#M:
XDW+:>[@@4EbBgBAT\FgXE33VbO7ZCW.a_?@O-dK6+^@IKV44Y=c^+GYK,W;E^Xe
b,V+N_fcc2MRYXT?7UPNJTW]PcP]T(egXJF_YegAODZ&P.bY-CYTZ9)&Q6HO6&^4
C?E:D^fX3@C]S#C82V)a4#8BK1QL7?8U@<-,,OQUE2W9ga)_BJ-<(PIX>V#gB]Z^
U:8g0(g/f3.9?1I]8/]Jb4@5G]C6S4A)3&cH)cU756?V.#K.g7]0D.8Z^4,MDL(6
?F><31]<[+M3AJF+7L0?#g_LW?IS]B4W6BO[Y+IABQW,AQV@-LFZEa=K7^XEO+HU
DWUP#]_<<OQ,FE1IT[J@(Da1d4WE\F8LE?JLAA0,#B<T2?6N<ggSI3C8D/2I@?ET
?UDBE.:B<gW(.ZRGf,bd(f&C>&bU;;@^ET=#1a<NXUVg_BR7cS1I1P4Z^<<AY>ZX
0a@]VI]2A3,Z@3/ANUA1BAI6<K>e>N0@ZbXe2@e9N6QV6K@T=-R#cGC^4C7HdB(3
=Td0Gc)c:CJ\eP=f8\V_M1VU:>=)f0D\__=(;SCW[2#\XLcA2A0P-)1Y]@A-_Q34
c@WfFFLB0E_H7b4)#a&_-Ea0NX6U)(GDF]IE3\&]BB:+,-E3V5_;,Ua^:8][eVQU
cAZ:V>?F<PCQ9MgI(ACRVe8FUV1<U]T19E3d\AK.7?==Af=O9d:aLQ26&93cME6D
::U?)RI7JPQ-[U>>V#HL=e15JDIT,d5;>XC@Nba_A,AC/M#@/5Ff@4\0[@-;);]R
4]#0NBH8YeVSMS:L>:&0M8WSSIcOE4B1W1[G?<N5WAY75P^<a7bPdTHA4#dUB+D6
F,->Q<CWT2@48):]G/EB3F(-[--<^R-65>,b:3>cgX&/eP/GGK_e2[JCX@T_5\.>
YPXMV#/H,0M:N3CXG<4-_MUP#bNCPRWAR;ZW<W#WBfW^6)L0N_C)LbFH;O&d8;1d
^E0HC[R8T18.gVFGKQ\:J=-V#_,X>:8)-\J;Y:;eOJCaZ733dZV]MT+^P1_5UH21
_X0DV](<HY0XNJXU@^,];G>VP.G6TE:IT\\cU:0:eU(#eYcK\J@K(dSE_KR5A1;a
U7dGeV;72HgD@[EO^9WHeeg@GPO0N+[<KBXTW0>U0983I\c>;59THMZ[>B^PK<Fd
L,GX1?XUcO,\dM^9>]W/.G&eF/g]?PPH2aG5\b3;B-c/_;9PH#H(4,E8/?N3?@CM
STVLD.+J=>^0<Z+8SNRcfL0.FPZ?cHVQZ+\2gN,RR9@@FIBLCL;7,WQ2=?eDM6)a
>1NOEX9DAF>U?7Z7E#77K3MI5dRKQI2.)WKMJ[F\C^a#cgadG4f5\\\#X2>a+AGg
FP]5(Id20_PebDXZCD^QXAIJ\S+3V)QHGITe5QA7MC)[D8SXfDHM7]8-FC/C0,&&
E8a>PU4E/F60eWVSL^O,V>AM@;G5O:[d>IOX7:dNN+K78G:3.<_b6d>-N\ObZeEa
#P5E2#X(9+2WVS=Q3W>Q#;.19@YED:6+EZT9T0cZKPZRd,K02[Nf2Rg(V/B2;(5c
XYg3/M6J=d^I2gec?5RLUN.0FJL[cPUMHJ40+79N86X,79T3?V8?<)L+e2gcC^/I
#9GB\JMfD8FaWf0@g1+VK;.&>g^H6FBed=GGN?24@1>76WH7Reg-cH>-V0BU@-ZQ
P?8[2>6,G:dH&&&;a])F(DK-M>VM9#@bEFPDC)H/FPNO,NI7E86,AFNgLd5VeFQ[
0\[2HKY6B:_Y&RX5CD[E(6E<2VFec<d;J6\^S05N^2fQBaSg?_K_ZLPe?52e=B(H
:GJ5bSd5:X)2OL4>gP+,CTMCA1?L5UWNPcXL=aU63Y_cSNP:T6SU>HE3-3O+\L>8
a\LVc7N9G\OAH5ZB7S218<@bWG3/-^[T;O\H[6aYI^VWRBYJf8Q-A8,+\+;LB\]L
-eXe<CWH/P:-Gc1</cVU;.H7@XCSI1X659g;A>7ZOM2=C#-2>\\R=2<MC&X5fGTN
IHOd@ee\1XC#M&Db?6:#]B[_6W?e3&&d^9>)U_#dWA;8I.WS0)_=a98;PTG+7<KN
DR02QW.Q,@+CL:E0]cQaL/6_cK[_e+aOad-f(.1H>#BO0FRfF1LY(XK#DHL=8VFd
N0@[[[1)GLJ5Ja8.L,FZBg]-RG8G&OU.I8R[[0O5Z)4RfJ0g4\M+f]Y]a/Q+R0-^
3Yg=dQ&daM:_VZJ:5.A;3e2[05>;+\?U^bV2PY5e9(K>TK<g3A9]83f^-Z+CB/O4
0J@cH.7NQMF2cYN2?@[_;Vd?V[1R&KAA6)fC>HCO#;P+1)ae.,[+Ne=,UC/OSA0G
NUD+[KN\e)K)ZPN]YHcIJQf_457&[ME[)O&&^H;2IGf:&3DW,IM=U\M(#+8EZfe9
EVFK2aR\19(Z&F:]2]R)>JU9=A>BZg;R3SS2L8LTP5N^3VU9#)&E4Od9.C+T4?LZ
FRZdOf]),+b-(Dg=DQ8MPPZE\J+OT9GM2^)R5d-B#6+Q/gL]0R^AaC-070Z5(T9a
\]VNO:O/P(&b:D5&X.B,d87A,J^FEb\T_S^.I1&d6gW23bP_3CE24-Z/Y,LHb2R]
6X2X?^NeE67dB=24IC[+I3-W@3NcLCX@FT+(;]c2R9;]O=Y?cD5_9K0b(7dbf(dd
.082,cH;Q9REU5:L9>S9(MOIV])J]abDNGWa=GP4[gQg<J.IY)OPbPcY:aXGg:O@
,eW.]/gN<K&IaKS-#^F&=WF(&dEUdP:.]KXcIER@gTA]0=gFgf<3:JLX]a:(P?2K
,WY\EDGb-K[e#5Sg)[d@,P:H#W[Y@fK3Kf<M)E]Ba:W,H#MA-90,g8;>VOR:9];D
Q]M:/Y466^>0;VKE,UG0\Uc^K1fA3D&ba.)bd3;&eV.f]8-I=,dJ(EEYI,,/0gNR
)eMEDc-00.T47[8_YDQ\CY[#]<IH^&@6e-Q8#+O&3a>JK^7SYE6K?UYc77DR_C)_
S[2+1XIbKHMcDb@5<HHV68<7I/dGLH=OCVc)J?SHBIDJ,c#(#?/Rf1Y-IOaSVT1A
OW0=d@.6f(/58PJU:ONO;W0YWQS#9WD?K42c^5#J<S/A-Ud6@)YUW-_<A7^I[U[7
BKbKBZQULTd;=PbTCdBeU1Z&CUbXd4(D11XUR,R(3(J)KfTDGW9IX=0>C@6A?UV:
:IEI@cY?:8:3#>ROfOeU5Q>VIR/cEW_<Pb/PRW<<GB43E;_La^aS\K;84.1:>F,A
YLF?00AJ8dA>W@AY,G?E7Q:B0B#M>C,WI#IM->5>X[R:^gNE4?dYT?2.Y^1B>HG0
5b+4D;)U/GRF[^:[+Lga9@\(<ZIaIZ8GNBX_TNMLC<Eg?e]&eT/K0AG/gKCM@dJE
Ra;g[aE&,-#?^=bEZQ3;c1-SO<VUIX,#Y1IJ,Me7.4g^+3-N1\NBV9TQD_#[5BQ=
L+&F8AJ5A.-W@]U,fZ3Efb7YY>LZTQ4(L6DPP8O(VS>>H<8:Df-#FJ1?GG8U(egO
)[;+>CG3PU>Y2LUe47#[H4;5cST8NNd(YI_Cg]70@RRbHI_M9SK7T-0eS=0(T<[=
#^]PRe.P=H_HS?FEd&3@eR.b:7,,Z\7>B;>7]N1[7(2Fe)0YYI4<7E_/PgA<,YVc
=.BZ8ZZI3EfXKc.^V12=QgT81P)7,>RRQ:?dGSN+QaF^I9(agPT&B8b+=<G\BPI9
0F6bM^R&5XYTM[K0]B0X(4TOa25A5EfY+-UXa83J3AXJb?&E[NQ]GUcY=S:@][dF
NQ3_-9AB>aNOK8(/cQ+QA\FM2[<)/\I^&2#[1g>WZ&V95N8Ve64>N_QVBO)B4?G6
M4TAQAR#]>.08GAb3JacCW[5(H=O1GW)c[#fQJGaN/J\E&>d>)5O-a=3QI5\ccg<
<IPO.]/gJ<90>EZXE<IBc@&WXfGDC1Q?D5@XLA7>+F@/QO?&7L/NfIFJ[8#+W[-+
OcNFfUJgFS^Xb?0Q1<[@UG^:FP8[PV-YJT^RW).EPC4YSaAT/GV4:]eTb2MZ2&(c
E>&-a>L#@e(V]5+@5(R?eIfGO&#BFaLF[B>CJ/IEg)Y=(:=dYVb/WUf>>2Vg[FHK
H(IBJfX:Yf&8cKVWBL\>;/c5H.^A7/PJ31>2DN:AHaJ;EHP&Wf4ASEFITa/+XV+>
,(JfEfGU8f=/WL#>1;<:=M3^ecMMCBLN>=;:(_F@,/FLXAM]0@dBPN&U6(#W9/67
g?R._@R:U(OVSS6a8;GF=FTK.E?X(_0E76M[UL[FFAJ)6d5bWcV]I4f2a-/gR:bS
-&7?E@&<>[1cISUEF.@#.<V/bKbEc[Ee/^H3FA+OKSfaAT-6GI.R+GVIa(\4V<&N
2b8>Xa6:f\8=QANdE&6Sc&6-MdA+;5831G(\V=.V?:PaR8_XTb;K@R1Me,:^:J;^
2G\/29g/JX-XJ((],;eXQA/Od#?Q1ABUN4H<.30..H;f-5MS\4+G5S)#6<g+eC4d
VU+e6Be1QA[<7H<\POF-?FZBEK3<[eFAOLS1=ZJ6Ef&?IbAL/+Z]A@>22,+>VTKE
MK3a]]b<(0L.f,0(,8;GZU9]<F&=EI(=U8De-BQH]MaXDR^,C/#3.HHc)SOB..\P
CT)1C[P4SHTJ[)YLdH)C:D=,5HAIVORLHHeHO=LZ5X&>QNb4(Q3&3^4Nc,27EgZg
fXA-E4J/D>cc^cL:QH>b.9YK^YgR8QZ(->R0]/]b@O;K[WRFBeW.]3GgK&399M/3
G/bY]61:013(G-dBEKD.Cae]UCSE(4^R][DgT</bM\ALT(-McKE]PF2c:f^/PU.g
B+6eZ)A<Y_4968M79CT0;0EI7&N&F->Ff).gWO4H>6_0H^@-@ROLcd?XU7-@BHTP
QgA^0DA[T_)X;Tca([aTeEEa8Xe^BdT2PbA8KR5Z#V^.&6YB/,U+,Zc2L@>-7e53
<^&Of0FI(X[?La2JA#-<=gc8CD?WPF3L--=g^.T0)ZSggcK_^ZV1g5=?0J9_2UY#
ec[7\6<=_^6;gAJ4aJ:=(YEA[)]#,1NYfb/WM6C?:9@?D>gBf@Y>:BgQ3:P&3T2.
7CA_(.KR<Gb?ZX;10TBbV[4C(7E6@Y:8FMGG0QVERb7Yb:+cPOFPF3<9([<5:Z>,
,?F<+K;&9,Yg&eO:1Y9^,(/I9g]FA[S#SK?R:W6;#E(K.T>JB-7_:KXeU+90<]7Z
g,XBcE=7WUb#(&1+_3J=?+7HFC,I,ef^+:+H_0KJ05U6#fSI@4D5#>_SeSF=N+1A
E5#4\:]O.(+G@7=YL59RG0K?XM,f2=F+9FJPc[;W9W)<7<6L>#gWR43LE9Y=<c3D
^b;-12G<#DTdNK#+SUS]X+cWXg7bL#G(dY4&W(K5@,9Y-;eE++PU3(V>&NNAA.T:
O2d)MT;>W7VF2X+6c1AeM2#gg);2g9FVI[Z>8#Le(&gRd+#-X1PTZI4Dbf85#Q?B
gd-<E6XdWFA/]@b/b9G&L9O9Y<.ZeF&EeXd+TVa[3#H_NPR&[DfUCf0-:MSdSF)b
BG#5S>EQC,<DDQ5F&_]Ye]P)[fE=-KcWKa[]CA:I5b@N=TDOBbRDLa_5aLMgF0O^
1T7Ba:=H1P(9J8CQGTH3:a]3bg++5>GD>^-?[IgYV_AK=[SO+27G1+Y/JHW4T\OS
F&1bY]9/Z^PQ_TO3GR@KH6Y&[<M<,W+02K5)87BGP1.0;_6Q;F;+P]?YZ99e4Mf+
9cc]L6P],BQeA-FWb)Vd(W?Oa<D+0gGCS@=^<P<#:ER5:U+UVf-LDHY#30XJKb2T
fN:F<<bcR]EQKeQ,Y<@LI[/>fd]4IaEE]S/932dg/6@a<2_R)H0=KH#VXW??-TRL
=1.<9)e08,fKTO7^+#eaB4490IR)EDe=U#B,K^]86g1A^H9NY#3eQE.KX@/8PP#S
S0BHTH2e^RIL?VVW6;L,,\YR1LLTK[-DVCS49LBO\G]1J++06(,Z8HG04UZDIXUP
08=;)_J36/f^1VBY6S)^,_+HYe879II=gU(W7ZH-O_b0I?BcPW0Ye\T(/P(KJaH6
_7gG,:QI)YYe7ZM;a;MU>.,?H-<A&R+:9f20N./4VQKLc:YJ?UE)2dZ54A6UWf;+
XSDa-)G;:R0.:B.V,L-\]fgT_Z154.I)+J&<QU_1NTI0a\31D5b8?<K+>#2f_Qf<
2M-HPZWDgUeP+#Z:.,f_M<b7B8998,Y&&X5#G<2>,=UAPWa4@56eQ?W3@+5+E]Wf
;3/;FI<G92fMUQe4eV.32(_ZS]&M;bceRE?00[5\X9a:+,Zba?K+I09P2.>C.gTS
B5_7<?HDP9K7Yf54]DX=N_B4;/2H-#gH8Z+be[;^-T_d#9FSEF79#7\fII>0DVQf
M1^Y@6.-B:/ER26M)0)5XL,)]KLU;),cJYYC@UYeI>a(f40/\Q?QF5P<:I4[;SW6
c@7(b/[f[:N)M[>)bS>FAV;VEF/Pb]Hf9H4XT[U=UJcaYL9@f;IEQ(&gaC[&WBQS
=U&0)MG3V_KB,TdBKaaJcOHIgWdQ&P[P+]]Q+02:_QPggOfDN4^EGB,-P_ST-0/Q
A^/J/Z(Q1>5R_QE/UP)aVYGf,3Ff5Y6afBa22Z..8Ug_:VM=^@_\B^4CfWPNEVZF
AJT8f,C/IZ<(c5-IKB5f0:EQP[b@9_(&]?cX6+S2[PD3-4PK04C2X6I_8aJ,TCd+
L/#+J]CW,HL2=7L;1aG31B&B<E]/#G>R#ecbNE7XCTX[.O+T06U:De_XScQ07+R2
)J_-._<7bTJOG:-5;32g^g33f+d>HP\5?[#RV;2e6b8efc-2C^,b_gJ_BeIDNBR?
J@eQWc=g&PaB0_c2-PK?<N[/JCbe7D]\OK0HXQBUbNHc>FK;^dgAK#OAEG/gAf+.
XZY,BcH?JGbNMR76RQ:MZWg[_&/[Q)\[\[)4Y>E)#]:4B@FaI^<f1)LWDMJ6=4JG
@]gR7I=OdMNUQe<1+T.X6^:5@QKa;C+M5Cc+-02.82BbC(NaTNYIe-XI7&5:\Oa>
C+>fM_8PQ&^P[OCDNR1L/UB@)\b6TeF4H1_ZJZPE_fY_7_ZQT2YY>K:=95d,CU@;
85GdVc[>MPDSZVVS[I<fEd[Ee>J3G_7Z9\Ag=O&eE0.6-M:)cZB\e4+^TS.2Wa)F
MLI<+0<9(;\.g,RB4ALU.QMYTJ.?7H;\EO8;-Q5K:B_C[3DJRM,?Haac9JCXW/\D
FFPDL2WV-/K?TI.DZ=#G:1,fPJ1\3_-:37gD7G)7SGTN6LX^f7:KFRPBWAfK1<5.
8XW?[f72+P<8K>;TL6e07EB1H4HUC@.NN_Mc]T+(T2d1DF&bRBE+ZD0(WUFUdJgY
CDaFQ-;PNWJ<,]<(dUYA>L;@G1../J.F[<NP7H,TG=aEJ;OYQUJS/N/WOXa3GMQ.
I>BNcQ)B5-:R_ac]+B)I=L^\LU[f7_VLdLF4XJ;LE;4gZ[8@Z0RJ>B>c1e/7NXC(
+VK?;?^a[>9C01GMBAA@IS6:7T9PTL?<,549W9M,b,6XM02@Cf3@WZJ#;C9+-^B3
&/.U/)L-+ND;.(Ie&1<N/]C75DM0.b<GKBC:fF+D[bVP]O6.I9>E\]5e+\F(d8.^
[;&:7AZ4YQT8K3_.T+=\2GXS@FH0MbRc-Y;]e2JGP^9,Y5&.?ERFOCO67N_0NWJH
c_5RGQ?9bbZec7eU<TTKQ<N(T343Ig,MI]E/PFgFQe(-F7IE:WbU;aF245KZ3K-8
e8[1UQF&?FL&AZ?8:-J?P8,7WU@V6@bF=\UI39Z=bJ4/DU@(fdgS(+4d6Z#^;KDb
\PE[0SPL2Rf&6/W.PeJRLA&PTR8]463^#I&/E83(4\(2<9dTF_XFF1gRK,:SCJ(5
H>55B8]ZB3RN/GG#_LL?PBa]5&W#RccA\ALdd7VDNJFO2-T[H>+?=S42a)&b#6CM
SYa?gA\PM8);&VXIegLf_4,#-OQ2R&FL>L/Ne)=;^7>LFWY8]AF^AK@4^ZO069IY
gJX_2&^==UQFPEaf48-7@/,YI&MG[KOMZLTE6X7HEG5e0O<4K/-F#eP(GKZ;U@2N
ND.dPXM\U8XEa9,]SZF<5?)[73,cZe+-RQB49UePa#d7DB+/eSRK+AGK^bW8QZSF
/a:CU;),BIfA[G_N?@,=L_\Y\QK,?N4^;P#;C/)AQ_(;;;F-C9ebT/d<IG^3AO,J
K;D,^Q>fG=)0W[f:XQG9?M<(7>1g(KA;7B>CbXRF333JVN@_B2b3g#^H8gff94+_
^H4\FZP.P(.Qd<\Db;?=NRFR3BEONHY/D1,T]TA)27=>T2;0b_N0-8d4S)FB>YQ:
?6?cD1T0Id&5X[P;H85b@,4&,(e-S9PY4;?AW01_VNdB?;/YQKK93?A=25=FgW]:
aN/5^5W6HG2bAO5U8Y3(X7^\+X5D1&-F\?YZ/O#)]JSTU0e)46KgN@#7GQ:2<YI:
1DZ=8BQK0aD<6ZIZ#LCBA/CC@+1C6dQ=E1MIFLbD_W[I5TN^\X8C[78a_BGO?<0T
KW=DN4>G/_a&9VC?[=^Re]]0IFJ?B/g3AB@eV80IME29&1[b6V^,9(24/DV^:0a/
3;-TQeOHWY^]>0a)S++a=N>E6OJVd1\&>(M7H/D,U]I8R/HJ7+a#[T&_F5RHbRRc
.>=MbGLf]_?XT_[9aC[<7XQWbQNc1)0-d/:LG,H<29Y5#(bf1I&A3.\_86LL.EJ:
)4]c&CFKZ6,FIRK@<@c]/g#Z]g9^;GRa+8\\3B3fP#.IAHO:e4e[>a>1?&6T\[#)
,?D7D+>MCN#:UD&B:IPIV\\6de7M>E0MYX5Q+YHE+RSU9:+.[)JM>RJ^A1,;EPIY
;,&S^.;\N9Kg1050dSBW+8ZA;]RS?I)6,fZLR@H7;B8a4bN\KSAFO/S6gS-^LW;4
0@N2Aae>C94e],_<f\<NR)\WH1NND5?f,Qe&_>7;5^-49LG[TF9IQ4^,>\MS?:-d
,J-UB8Y1@c,T3aY)Jg/fXL2;SEK84-3N<_0YCMN5:f:]=4[9bdZe@.d;17F^,_(f
dISBc-G(9M.E9UB:LC^\2ZKEY_bHS3F,_PDEb?W23S.;3U)Cb1^MT/J+8N+>(.W]
9DZ\7N&Pa;BIaV9J<#eMXf(a3/&X\(24T4QXe3LagL6PAV(X2C8X)GK=<AOK?],(
TW4+W<;PE\8DEQR>RXQ>+&U&GQ7IN8dF5f(@a#E0K;?7UMH+R<f/U2Wg8A0gT5;0
fD5NdOf#M@ZBSVWOK&NI#fN0WC7+Z)URTE?A6B,M[P2Of3aP(NE_NUF-=D0C:&F9
?<R\RPCOGW/;>AT_=gST#H([A3&E5@O:W3dEI&++YS4?ed7f:.:&A5>_2gXb&HKH
D4)J(&R,SK4D=?g)^,M[>^ZJ_A(LXY=,CER9[1V5Y7-I)fJY.^^OFdU&[8e<8Cf^
a494REI#Y9C@E+?DA2-YbfE.a<4BK<U6[;(&S;3[Xdg@Z3.b:]acd@5YB;)Be(B8
Y-)dE?5K\DdS[J((gHdagN:K+,2SV)#-&dZ;N+7F];U0CbPA(,gK)_\SKB:[g9F1
E5^7MLGcB-^C&&C6+2F#W1WB[W?HECOT6T)/c(#<bDU_3Y>Y#9gY4YDNDWSUbgcX
)IH9Z5:<OJ4+@SYa/Z93Q=7YX4aDE&C2_C=IL+ZD6b?-A2;TGa(S[G\6HYJ8aFV4
\1SKEZL1\ZN<H&#5;HT(Gff8528Q66)H7BB9BR7e+EFgTV=<db3@_5(_Zcd=FS7J
OeRf94]I(<\H+6<O(4&S(I7c(617J0?-+U;0dXUJ;AHT(OINV@QOWED?&L\f\;ZM
3?@IXgZ/H@WXJA;K>_&)@4C[SN]+EOB\2^-@1^4P6<P[&f=5.-TDR.>GD8XLO\Y@
e,\]:NF=<RM=5SOSRJ1+T?J5_E=Mc6=432&DUB[RDQSN5.\ICbBR-<b2_2bU?a77
WZS4WMGMPD-Q\[YB9[0<;ED(Da+OM&)6(B]MR7NTCG\e52+Q2+c9We4=XdJ86CI1
SDPN874NQ+]F#NcY4..7c1X7.HS)g3.1@URDB?Ed:0V=#PAH[6K(^/3[C6U@(]Wf
G7HFS_\bQ:Ua(O[]56_K(RCB-[#=>-GPV\7G,[,(=dNN.A7e^(XB0D9USP8#R,dN
EbA8#G&9d8F5-,P:+=#:J@?gGQ^C,NFge?_D<b_.P<bK6:e-b<6F:BM,#6ePX)Ff
GX;[HS3RPSaN)K=)GI5=#/&)GNd^5c&N7:]]a\F6581--XHbfW(\^ZK(DOZ)5H2K
>P=d.-RS:&\BI]35>/->SF@;+=VUL9(?#06C:E\=U^c^B=(02Y,(EAEc[S8Z8bUC
3==K/Ve;_^JASF+X)RTdaOY;.C4CYDN4(I/;RP\=+QQ@<?G5&@OIQH0QD>S/bb<S
3+&XPR3cgP2)5TZfNLYaK(JX/LQS):2D/+L5GW4@XR<D#Ub(JL8f:LB4GDG@E30F
68+\CHXH9:_>YT8SVXK0G_:Q)/IT?P@:LYM.OdaMBbO6SE[.YK)K#=c8/#c(KSYO
-ff.0OCIbNR1&F<VfOSI9a:KJ8Ua[L,Q81A5NE#XW5A,T)[QBB7TU:E:3Y,HSJ5A
?+3]#[^XUBDB/HO+AEX#K3)ND(/&/GUL5]KVg31)&.6WQ_GQ/RIXG>O6X0V/-S&@
LT;Z<X5+70]3eDK,M3V@TI5ad0I<43bK5K@eZ5+g91(CB9dIK_Zfc&d745\gc5Lc
&<4K-Hb1F/_#B)9T]^f<XG=>^O_A2)O>18P04DRU;Z\H/d&6b<@STdc<KeN=,+ZL
0EVRY^bGJY,3O=V=<b]d_EWRVEC^YC89X#[?B.8KBFMQ:2D>I.P-R4M:LY;:G-G[
.]N;=JKbQEU+FE#D0b/Cc/c&.A8>=M)VGY:;?7>6GHf/<RKYU;A#A(+71<PTJ>e-
#?U#@bd_].,c3^,YZ76,7f#1:-FVefF07[/FJLO=U3+d41[8fV)a8PGZ9W6ba.Z#
d,6RM2XZ?QfNgc[6<c1V\)+:6U/?VK?N)\0cEf<,E<Z1:EMZgZJCc>[6Q[EgYUO<
VeMA1A14LFEIPQSH>B5G^VN,&M@4/3]&G@(f:@6BX0HWDIF[fC9V_G<c)N7^MK0D
VY7K^\c=YZSR<D,3CXE#3Rg2&^CW=6]gHa\\:MBP6R#+@:RNHW::<+=;OX)?a3g-
aK?6A306Mg[1He>DEP/(&U1X#Pb?G.5>(bH,JRgNf>\7X^=HI.R[<11@@S4-.:YL
MZJQ1Ze&,52<:0W?H<B+bUPK+>F8UTOPU[H,[?@;]WDOCR;C3>,/>G.<[bN[,I;f
-2#A<T(A?<AEVeeL)C8PI#c79?J-N@F0:$
`endprotected
endmodule



