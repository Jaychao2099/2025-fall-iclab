//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
bNLlZfuVqizS4uhMsx2n/kaD85sq++L6SyXkV3EhNZjGjJ8fu2FNSmFLWrvPo5CO
Q9+s80UgJP+h7BDcy10oXiUJk2XU8d4q7BtWXGkJJIUQ8iuH0H/wM/dUi3t/6k49
0aQduLQPrrUKXqbZv31pqndirrnYfim7jIJgHDaj34rPlIpKE8Hc31VSZL0I32bt
TZQ9kjjqV6Vr4vkjiKO9Z/1BxVIF2hdnMse5hY5TsS1Gkpl8h45+6I9k0ZDg8SnU
CvDlUf0EoI+F++i+F9LiRaJjroS7IFIBEsIl6atFGN1yGac/Re04ML3KbO1Zibg+
MZAaMv86jvKdwc63FrkBIg==
//pragma protect end_key_block
//pragma protect digest_block
PpLW2T0kzkEl5ZZeFWXnXIKM4lw=
//pragma protect end_digest_block
//pragma protect data_block
CK+ot3DQqdXP+OeGaURM93HvslJj01LDdxv0hYhpldP6ihPEGEQLr6ZS4/6pErzB
eBI2RVypPROYoYshqfYWnoo7UhXoQNcsIFI3b621tXiaQ9GDTMFdRmuzs297XeNN
kvyvmdvTe3XC8pvxwzDAQ07Z+l4AjKnNy8AEinteqo1L529o6rDqLo512Ebbfzi9
H/30F2xCh4rC7y2svwtyopHL2Og40qAjzBr2t8E+E1+wXqrXSOyJ9v/vThYchGoC
WBc4E3ptbS7kU3RXJgN7oFmC6k77qNU5007mzHjSrj+VRkQ1JJtPkkdntNE7TQV5
6WKEeTA3uSeh21TeS5IhoHzURR+kjYc0YnHnyrP6ozGA++Ek2RI67alyZhRDnj3T
ZbBiQlqkRnPf970Yl5/LF4E0r4o6RItH7PMH8vhKU7wfuloGRbk72U4JtkRMeQLK
r0A63aCbJ7NtoHkTRQo3z7VclHdz2kfkOhUA03TQ3Pai7BwUjCOoSGdnb3F4Lqri
rYG7DlNcJX5CysDxM1aCrr5/gp7f8pX1n9WN1gBYMpqPmHV6Dz+a3YzarEeUJHL4
6R3GK/qvlcukCbfeJv7WdKnhXqegnXLAm1DM9Os8cqZKwd4FXr0SMn6xSYkssTt4
kwrBzl8nSvuIB0XvGBvb6PE2nH9HNVbdcuXcOHP0H3VJupnxdUACO3ItGA73AWqZ
pKXVcDfZHjDqZvvqytNtU5kQLJpbCXod2d2aYSXIPl7BqTAaqBUvLEZHnEWoK1X4
y57TnYNB+OPodcruoU3DuvVNs4t1wAGhrzNXKO+gtgLb5Ty7GweRdKsc3g8jfpuA
XL9Nx2+aeydKd23qaZadVsyhbYkv2HbSFqsTHWIUPQmKwAqnjG7zJ7RNAzlzSWe3
0Neu4IlYCzm9L2FgcDtj1lEXJTHs222HdvtQduuB+STxF5UjbBXgT8XFkkPoi/HA
cuR4CYzxRvH1GJwhPD1yL++OXPqTKonB2T3fJlhF/YC420Ro9pw1cPMz6n7k0B9A
mak/fzLYHS7zfHnu5LIuWgb0i6JAPVCmwvfJGOyUfStGwnS29YttYRtITGJC0zWt
K7nOVOSW3sSCS+32Rk/nuEhvbNyPnx9hy0iANaTbHHp+Z+Xh6IvVEkdbKJUekqdI
hLdpaGd9JQuVZP9LaxRIiX3v8jVYN20WQK919A4ctcg+kT6DPaHoEPhn1xG5xYH4
SQEz1YzR2+wHNi7Yz+QwLU1kiWPvwEoyowlPVU0s/9eoHD1vP4k725JjZ82eK/aj
qm/T9UI74VCbeoWZ0lOWXemZv0cmGIQsiXnCqtz5RGQu35i/nvdBCTnyNSYmWyKv
o0A1OFwvmimJP77C3qBoitEww465ibQ+4lrPsFCVYm+bpsIZ0/7HOgjfV52pV/+t
e+6d992IAJZ6WERYC8bwRBnAixgDLHIZzsUlXdPumsyGAwcOLSdtoIS0ucqKswEx
4so/CgV+KsxOHBlCT5oj4DgWnV4Ft01BNqdAduMKiZsucbQuHp5ADgGJcA/RISVf
J3yR6/5jlIweo3nSuCBFqZeVI6srQyagRUYvWrdbsmTzk3b7f5IiEbr94/dAuKoy
Y5vwRPoe6pHB2CXb7ULUksRycNf45qEIWqlajZZs6fbMtDC+Efpcp32Db7C2b1kc
F+xeZgkhn8bzwIyY4gFBZvpcdICxME66CJmo8gJojQxjJJ83VbCkPKFS5J0v3wdt
QMoxxgZL+dn0EJ3IYUYcZCRSHy+1RQfSvJk/Hp+42H2aBNuPnbgpwRfbvqSNlSub
ePXjZ0PM7NmnokHiUMVDJMNVoOcEawHcXx8v1VFaLFqkxC+xq1QLz4aCp+0xjpal
wltSWJz7GBjCX10erGBhLNdO/KODEmf7X567ZzGigs8PWgc2aHRMssYcFQwyQEEy
UQAUnZj2EGtZUECPGQVrvGS0k8GkCR/WyzEHXem1yTY4L5OCy9qVHFJj8w6bErHj
nF1RkS66WDptlV+bSK1z4WN0PnjotVVa6BT3U8mdYv7ANglW9ORhN+wO28tOVuZT
OqAPlq0RTsNpULMiuIRpSTvoIEcvW1nUIvNdq5nOW5j0ayN4Sr1NpNI4jFjNMwd2
LHMlbCqbabUDUO7CZnTxqiG4P5YbDy/bh+PaxIAbjL0j0OPfrqiEDiOZQVDu5hW+
Fp+HFRtXIJnayF+ahZFA4sNIwfkRRsP9dJ8jrd836T/ACp/fokCKer+pA3zeTWb2
HCBiFrNsjTdgActfofgB3G2bS1VVn2Ml73OL4eioGfKPE4eJt4iOHF1Ni8dhIy3z
UrYiv5tJwKFJDHZ8CyN3we6G1vATnY0wTdkOiYnq2LkCTPvxhGag2POtSU6FQCzE
jqnOATk8HeGG83aQFfCSwch1BwdI1ESzf6z/RVXEkoqymrZqH1XifqaU7tH3Rclg
8karDdZhtbSA1GsT3hS5/UvrcGx7pA+Np1iCdUuap8vpphOXkZy6yLxyqXiePRp5
arnK/k7iySIhzzxxtoWjLJB3Gyvbel5X49ocoiW1//KJdXhhh/PyC5PEL3K0AhPB
GxyPtD8H0P0Wap0fMLSuCRCvfhMUN/M3vmMHw3BVXco1JCVVq64JLT2UxYHdQ3/Q
4dtmlgm28EdnSu7R+cfbJDjlxQ1jWsUPkWcgofQfW4dAmzbTScnQDlwwg0fsTSPi
5YjpR/PzN5qYDOtieq9frf+8hn8ztMD+iydKtXOJhQo+bLGESRx15rfW9DUdHttM
Z7xQORGWUA2glXIBRR6fZDpcNYcstfuhTN5+vd/oNC4BI0gyq/NQR0U6TF2EJSJ1
Dl/OOZC4egHE34t6O4aSBM2xggaob0NTTHnxdAm08DDdHF+HzYbgTOcVFXRxVxJz
2HHL0YUE3USja6z8KOYm0TnOBaOrZOspzh2zSAT9plmcfotrRfp/XAXVOr4P/+iK
5S/wwciAkWcRFVAxz5OHc1M9yK0a8BixOFPbxarKlqXQamC3DN/DFj6dwuozBT/1
kK0zVAIKBYEqU0CwhaYKvT6hyTxEiUL399YxWcRnlrNpDjx01bnu0h7RDsCnPD1S
IKDMDmqzBKjXjVMcd+OrQvwltYBeP5WYmeGyP687SjvDCJFzQIU79EXCNXkTrKBa
ZSWTGeBXf3E3tuFU0WxvP6wTSx3eJTr5idHGQVyy2k2yXvMBMQ0WdUPaFdy4VuyO
B/EsOcyHkLFclu0t7qlwITZxGiElAo37+HzGOWEpFfe2rXOgiKrzZZLJLlemGFYD
wPsNgt5rnfpE3WLluSc0MFYF/dYfbzj991U5ioEMn+ccLvswwfgxoUn6PikYKW8S
g1kotLrMEiD9pvC8h2hiUUTIlmXT3gTRgCl6KIclnLMogoCLeam5Ov7gZrp4G4rb
QnjIOYHsryA4B8jJG4sP9ckl6anvYHgoISt1CvUf4fjoj+6EOsACx+HPqYxMv8f4
x6+Kt3OAF2VI5UTFu1DHzMQsLh9ua+UGCeCT8winxbnkpO2kYWrXHhkEGshLkpVx
UPmM3jjgUhLzjq1wA7raT1PUns6uYRo9uKHvlaIKiydrQiAEd3PoqPb4H3fSErpQ
skBTNDexAWEJfZO2tURiZWkwtpcEYhEnr0V6FFTRiFfulF4MrXaPDbibxLeyZgkt
P9S5ba4Rhxy9e++0qwar/o3tMDczje0RBKAXfF7gQCTUoJYp6Xoxg5V+8PQXBSv8
BkLQSgzJjb123E2QGY/1J6LQrn33BBmT669zNxUBwQRkt0NM8qsT/tEGh4CNQ68E
Fii4HqbjpS/kVBFTgBKup3hN+kz5fqvOklryuEuo61hlbi48Jkrcwk8RzUGe4yDD
QBlaV6OJsSN+HyomMY5YjsWIHEFXFhu5ZzDILecB5F7FsB219uD2N7EuqWme7HaC
DuyKr3iG6MXau4iXsohTiosXOXUdrJy1WWHeuz2obFzLpbSjQVAEUXmy40jPPqaa
kkcgCDZDifS5Cz8mTYxm8VeKQFmKZRmKl12IUSxzRlOLm6io6HluF8DyjoUUg9dp
/n0KCc4d4cAhMTmfzgJUWLMj4BF9U62XHw9eJ7AIisZZ5vpRGJKSeUysQ0jXAcvL
Eys9R1jYUTYVpAPi17ygbb5abMlzm14zJlZVPUASZuXLN27T64jXb6rRsc+nXh7C
gzgy5O1ONYjP1jlAkg6w0rmv7uz9/350nSMtHAx+tWO2skcgTy05V5Cd5GacS+nN
6TMpQtoQYC8iWA+zT5AFKHS5+om+bTuzf2ik0kaAUh7v34otpK8gfIkrb/01aDH4
GxMxd1ceTTPtO71uULQEJ/dg2o+yhnz8FBAhXm/l+j304rmTDSkVgd+igm1vtCqZ
vNqfEVUc8Sw7RWI7jxdSCUqaLNYjra0X55ShI6IG5ikl50wzwSGjgloGufYLw2eS
aBsW1gg3PrXrAwyrDf+U3si9t3QFsHZ5mDKnpv1T4r5ESqlF1YyGfy408D1D0AYj
EOHpqd1FUVnJIhEy1EIaefQd+n8yY4JizfOwKBSaSVGoIlQ00D/7IshHe2jg0MEx
oYUVdLThT0941pR6kELOWUE/jliZNTEdA0X0ikhkC61jFu9uQc59tP/Ljcesz8c3
nppi4j6oEv24P6b6DguwC6GcYHJA85NSQavalFOUDViySagpoyqpYbZv+Ix6KLNw
59+AG4JMmoOjaNzrniVweXcZhaj3hTTdfhw6ps4sg29vHGLHHkM89ng1esolA87I
zKFLsaaRRekt2bHXAYz8ylYMM0oBM/DDkHN2PD+0AEgXYsw2/twEZtySL2c8j+jA
/+lrjXxbSOmfrq+F81rzMyCThYnersV11eGJGGTQxwmNhjq0aMgNUIKRR4rrW1LT
pfIf7ZZE1lVaUcPSNoKogX3IayxDpqk0jwMVmX1bp1sVEEdWfn8WO6LlQ+KJZJiY
YMeisL5sh828hhrQaluLJsQmQYzIFwdDXDOdxYshqNPVw+bggKkaLnLmzxye9K50
lI59T2cDQSt8a7Mr0qlh7tzaBK5mjm0dMVkI+6q1qU89ptrs026i9j9822gFXTWT
5aqB6Ox/Wv/BlFqlO5BqhAy12c1L4OT06F98ZHBvR4kFECKopdUOMM4fnYbRMqmr
8w9/TcTZgxq9S4bbPdls0kloKxQnlTNsVS4mj6kj3RPhGYoxkLhCWpbEZITai/Sy
O3+iOl58u5AomaOdsU7iHijJpkgDMslL30vwICJGhfEmqg3tAB1cKd343w9aofLM
xLgw2Zb8+KFSflVzeShzElNOb5bXpoC9KmE0sRvrkrt/qFcPFam1+bymKJ2gp+4g
QJ0mLBcXL4JGha9MVJaoLhYJPRz25yplMH2zSK3t+TrVSCAoUnrI7VISht0q8owp
TJNqZkA9wZgE8ZDW/OMl1Q0SqhttUAgRlx2RfRnNFneL3Qz/0IH2hlQNMRpdwW4j
WafCLIFfC1ukOIRmq9H7XRUISUto7QKgHkogHoc80tA06lCF9VU1N9BVfaVVtK8+
XNGjyOuNItpWul589VvdOGfTx/39oPp+N78/VinFS2oTobx0hpD5HUCnSdVF8KXw
HBkn91OrR3FuoZ2O2qqnnbGQ5AYwl9a7AjMVsIlEGffQqiCuBOWiOqI5uKQLl2Ab
mbbl50kH175UT5InG5573Ibhf5ZPdv2wYYPObLUIpfwl3o4n1rGKaUZOCthUR9xZ
UVCCLNtRFw2ALrIxYklh2lyZA4HO/Uecp+N/YIewbOhZEl1jiE8qR6e/kA30O9Oh
rn1bIfExVAemd1IYApJ1ik00asvAfSCQabVWXTnE+ln/cXe/Wor4iKSvGj9wPKda
uHmVjyjODQN0WFdmwj4qdBvMlohLAjNQfT2al7HwBy6ubzP/jGBaNu8S4Iz/g2bg
uNz7+cx4Bh2eS2vtIufckZFaka+b/A1lbtw9HBY7GIRqXkWugb2OCrgXisVppCPD
jHQjRtt+fZXUWENi2tFG928YBfpmeMZfqMg8WXa7Vz8a5WXI2NG0iZrcH2oGoNNv
nk0lEZ97XN65MTVcujIBwd1ymF3rVLxfrp0Xxvd0BiwACoqt2aWFGq++OtmDMF5z
rD623ox0Cf8jtTXqeIpDRbt9KhO371zYqM+irfADIe9nCkVQp1On4+OohTouR+Qh
mpRkiGQu9f8L0Pq/jGIZGthjTyCMGUPM/KWsdEiJDOose8nQjUPu7HIM4qbgTGKI
bEA4qtE7mZKOoofjJ639lBPFVl2H/ENqt1KZiN8vVy3aZoZ9TjylioxKgg1Dc8Tz
6NLN9Ced3ZjkfdVplZoPIzi57KiuGcN5xTFa0U15KT91mVoNx1c0ECWfQ/GhC+4V
j0HLduwJedZd1MzCBTGA9req79vlWIKrnGRPi1uOGyofvrzhNu0Q4Pj2/o4g6M9v
CJR9LD2XMWJlD7pVo/q0SVm0qHnVcZHHESnmhjshWq84c2pByRhXtRguPRm8or+3
o3Xw57l1UVAoeYOR44koWnr+sXZMC+a2Y5dOEO6NoO9d9OVCHMZVm1a97fU28cvL
EXXYlfzXQvy+6VwujJunW2MCH6gtgxYoGH117RnIIbtR0Y/q0cvfjxiRVVfGAjna
mYfeEP1fdWvzvxui1zUBw0pSk0evQ+jYSmjZptdhVD8AHUGRhsOLP8LMv8J1/dcZ
XFQuSYEDcas1lUdTVbY2wBly+EnskxcNNQ07ZGoeHdGEEjqADa7rxg2sKz9tBbXc
sNF7Sep4S09kkD/6MYuYxuU+Y0NLNAbLp7t57UwLHMcRcj1QUc9+nzJCnG49av6v
1mIC9M7SV4t+dB29j0JM5rwuH48zav7nd7S/iXWtuTJVob3jdjfWz4peeox2oLtR
5bjSWUi45fO2pcPeigPeO8Pm5kSyXkwPzn9Kk9Id3k6a9k8IT5+IGkKfLJLLCfhb
nYDxbHyOQrJzzEoA3JXSjA4zP7tECOfQKaCdyyYBRn86YcKYzMmRe0mIyt+MnDMr
EwNvxc5oqPyVTwW2hjVfrVEjG1xyty88znQNlNJwsdR6SuXqrwp+3v+0czZPmtcs
0ozLMUYb/QyZ/d6BXCmpG+1cHfhkYBN80VEKfuxrCdksxoWqP3KV/7Vx7UBRjCTR
GfVBKrGYS/JPXcaG71ASLGktpurXR80omkNVxRvZ90oOwt8V79jhN3VktIcf2Cd0
7HzfEilUJhg8Q+Tg5Zm/aUXLil1xROHt2LcqPMuYS75fImFTDENV0sV6xf6ZezAn
TbcsBIZBVDQ/4MNn60t1OHOxo1L2WRKQ9YvMRCMo++dIL8BEj2k2hUNaoPCxa2z3
u3gvmpi8thtrQJW7fVKiRnySFTcZZ1wGyrRKLzGvhOsgGQU9YPS2lkAfx0BqSDus
dlnqXVniU11ByHxleIvUyba9q2R2/EoXh9CbaOXRGZVShjpAdRNMxm/iBWgeFB3s
vNseOu29MqLtY0IFcaGglWQ7zvYwQMid0wFODWYNu/r3KBu5k8iVAPcDlix3i7ZM
1WlPt+I+7dFInYVUG1c1vFLOwQ5ea7mP+iDjPsKykR7YH9B7UUos9mL7vkr8xtiA
pdbNUfAOEgA3MBX3661cz4dBRRap+cV4cLZ2AwKNT1CEhg88Ur8Ecb5YbHS6E8gi
u4pNtsCwUtMDu1LkjnAIJNDp8SGnPhDwpS1InwK3R4ckvLRCNkI/Pn9qo8Il4PoN
xr6WI8jcOCYuECf4iwaKMGXVrn7opvHT0C37aFfYIH6JVZRoWTJNdxEztI/1Vgxv
PovHlNXWDgjUv7hDZyFGOlt3iaiVWCXGeVdq3KIQr8qgOq3H7Bp1AeZMsiH1eFB0
m8MD8+jrt1AzIIT9rlqHFuDdVe149QJFZ7nhghd5jOlunDW8eQ+vQXH5TVfzTujl
hLBdMASD0a68Ckb9NfwdQMAhazwaTzJ0RotNzrODTiRIVFw7R4H5AF9sNZpw+kw1
TgOVmD7FL0jrXyV+O4b3ARSgSzI9dvjMrv29nc3Bx/BqZtgxuay2M+CQRZwViAsp
TBrd0GUhWr7YNUDGShBNJLXI4l1o0KZUDUm8eiIiEHRNd5Re90SeyKXOkyHdgB7M
xYpHOhkD1haqodRLFMbDwVMAG22LGlqv513dLoaOCyvefym5oJS+/dlA3APLt423
m99pbFWs08IoeEBhObzkLVDJR1wHsKKh3kgLdI2H05KxU1g0h9XnIm02sndpjIaA
NWfwePSo6OQw6/J20iT8tZeFCyQ0Q+8v+cnxANQUlnUnOK9uehnmzSASK7i1Xqm2
mSf5GLjLUiOsI7VOZgAd5pFQjBhr8uogR4bDRmevCFYzH905RMVoe9cca7KQFBni
Ox165MxFF8AxQvv89FR4ab2AXDadi3CESGzY1m0tTMY0lNOWza+RTCMyEDD/3MEx
k0gF0CnMVE3iLVbsL94bUohBBov6Ql68rxpM/0KM+jpFcTak72t30Y+JfksPDdA9
wge/9txJq6V2hrOiqKWTps3h8Qq4Xc70Siw9O3ebI34ZwnUQ45WLPQ3B7Mh9QNCy
w/izKtHYAZy1y/FVMjXkLOHVyK6LRKYTbKF7cSTsa5cXqjEsi2hvC740uUJFEVPV
wIkUCpbWVB88ctX6TUnP0n2mCQJ4sETPXnb32uPr13BrxYN0ScthoVVl6tWUxJMb
GlH96cpQ7lWyHRTNQ1OR9SnUh6+GMtROlvxpRsPSqcDuhHIoxgSoYj0ifzKw+iH6
a13IFlJDJt8yktH7a/A1yvUBBdm1PRyMvC1yyhGVSmwXVfLg93+NGYfdsgvA4ecs
EPbfQrxgUK052XWTUzA2y2GT63CkFc9z58zKnEvZ2W7MYF7RvWxvIEWmFYFXXSmR
j/J5+f4HMHa2lZjKQ0sJk2hc2ERJNFr2hmOPqUzAFipoPeRil4G8bCZ4shvr7N4M
g+H8p/iSnX3OKUQjExVAXbEN3fe+VpCkb7NM8u60H0URvVrqLiqvaHL9amWLTO4M
gsm/pOZs6kkJzT+mIbSs5rH78PNzd6ocjVYLTIlF8kyLzs+Gs4Gxg6wF6urPGImd
lttLazk5Y/KaLYHgGLHE+yoY5EWGeEfLDPWD7NpLQQK81H74AI23oObwp1c3anvQ
ZJ9YCF4TklMj5mHc1bt1uCzlNUv45hmTtAEasKQ9t0rxL+WblExMl/XpY3m+aAU0
AFYccyviTiLE/miLDfT0iUCWeHwnP3F3Vi97eSiCKV/fYngouB322vly3dCs3nl6
cIBW/tA+WGnWG9Vft2FJxjm9K+xIBS+NZTUdBea5P11zTpQzafglTsozTpb7Z+OL
UQq2xSJLrcTB1xQ+jt1+BYPKfQi3ZYJNB04cQNVPmj8Qo19WobBIugNzsvIZwdKJ
prOaP1UK19I2rwMx2Xi0/SMSCbFu7gKerR64CyyX5Iz0T7Dc0651TQD0S360auuj
ezI+BIHkILOmfhmr4eC2ojkB90rPzir192kZZGGFIGEg08poafboM8e8hccpkCIS
+dx1yRp1A9eGWHFwn9Hp4nJETilHWm8jwMMAB3eBhPon/rRtBEqmYJfvU80VslVt
CEspQq7AEf5tFvwFA3i8ihX8ejd8dngdduqJKKRkzCRvGuCV+Q4ndMk7P1c/rCTt
x/fb5PgX0wxpWk8Lszsb5UIW8tE0MpT3AD2B96YOwOmdMCDFfThQEqoGPDAe8xq3
5w81BSEsmHvV9CKFafoX0OA2JskAl8ZcTwc4AqFbrksWKHaWspwdI7ZpXjy7ecLm
EdxWdRGZ0XoBdYWH5MUrNkGyL8xw/oRQLtya4sBUVm9LAdKBtVmTvwu8T+NAciYX
gPG9FV7RhEAhtHDyYLPaqn7Yl+HqmEC/ml94QVNa4VO5KB3011TeNM3s8z6FT9dE
OfYAni/sWWnLoLMBIcK5mh5TCXxxVTpC+oSyAssSwK35VUc8BpZOtTacpKu1khgr
nAxlUfJLFCa665to/GcoxQ4YxM6ipiuxEmKCkH4aLdQ2utVxVNjbR0ZBklZHLGdZ
L+SWG4hqQ59A8oSLcFUM17/7I8v6gXmfCCSrn7fiPHFyf0ODCGdk49W64nimgecb
nAFqYpdR5wsnecwTEqbfOTWm17pmveSqYIYuwQTm1BoweV+Y3Z6NN7EHlafFKdKX
gwskaVJo7qveF3K8/G02XD5e0BfxDYyV3OZEE2zxkgixzELPawaMf6XTUOi6D2Pv
p2NmVer8L3UkegS4TGNktaBhKu+TP3lihrQTzydPwhARO3K8QqFbwWGv8/2ZIT1L
RpkS7eQk4PBSV2sOZO6nw6032WRFhWPnMh1iTqaNIFKQ1aFk2UKqbF+QTowewjmy
ui8OqA2/OFUGYzZB4iyIoTd4U01/B1sRlYhguG21Dq8vNejU6sUsk+rXxom3tYhw
c31MwGWq5Yjlnnnafp3hFD97F6VdpEyDMalIC8jrXMK5+R8fkQUMmdEZoCfMqhaG
zaSlurb488pTlSGOkuD0pdBkEYsnjkc/gQsP3zXLwdvjfUWsdYOPfwypeZSdO0Xl
EJf0R4qqKX/yc1KQFWZeqUrQa+fGbFEDwn/PtNJuLZ4P844WbDxSXSf+YoJxYbxg
fQP1DJzl+aLBu8RBfKSUrobiFmkKNOu7l9V5kyJyGLEfjx9+3EoneQ/jn1nOxu8X
T9+sIqMNxJ0Ee2HRp/IimQ06QCnlAueuoFZpzShUcbFrhZewNium7LvSvt15rdo/
hREOs+qCvVFyBjCxpH+Es9Aw4xJ6v9ELefLo7cREcj9hk4fCzCjQoZQaGHANcDAs
nGK477afpreblp84xLROrAS6S3GVPA+tNe4Kwqjm08ts26aNWlKL3UWZeE2kh37s
AS4NLi8cXfVrPqKxsUhkaLJN8FqNwt2lxGNnQfpi2ZojGd2GRHrkRjRhZfi4AMB1
P2uSd7Butr1EC21z69COxAxtqBvZeAMYAYUEuI3GeaS94dKy4t2ufI3yc3NeOt/E
2qnTWADx8EpaMtV6tuZQZwXjSXZyxbUPxwhUsuk+3DPKTxakJhG0Z3h1JSJs3l++
Yg8K7KVISbBrvGdN/s5LhJXu1qNoX43XeEfV9Y28wkngUt+2harNVRkCaYK/ERPY
MwXXpLTmrNAvehRHmdz5K0JzYLUWLI7g91R0oFQzOeGmttAjXa2shnNKGDhI+8VD
QBOuTqdsCE4DrkPn9caIrNdb/NVr2RGfOtZUSeb+NlTBHPI0btMo9zSO8XMN2oeR
9zPA73+rw653jOsM77iQMR8mvpFWXYnI1qo9bKe7J5rO3vEhVwA/ZlQuakMjsK5C
oqvTXl7QvirjPE4kaT3yKUWN76LK4BUnjJcAp1dAjyD3TgDnLWKMt/Wtcg0k7q5x
2a9QYyfkPz1Y9ApcL45h2V4nWqJc/xWbTT3wB4zCl/Jj0j06CQqN1AlTHasOiSAG
g8M29fkQrALB6kowuBPAhvr/UOXnwHcVziJTZUTDL2yz2QuOXUK+BuzjTUpuqtt4
NraVXIMg2WY+5lsPn9aWqQI6cwMtt1qNeyQ3lTh94bm5BbyEV2L4luT7ES3MoW2X
uUVhxOyXX8zefqPc3s5n6TRQQ6Zgf1ZZ/BMPk9iTc0f3125YhPEvBMZ6Is8Ew+sM
FRuxKCDYOND66ZPYgKTEJK21KNJkKK4qhDs7hLUrLeLmO9E4k+ogo+5NV3Z3QyNF
FGeaQw0T7Hvu7sj0K7b1sh97x+clRd2EBbcW5y0Fg/druomKiB3+HiIUyVLOLbnO
UHdfHvB/YoTmV/+7n4n6+bp6dYxEdiJCDKlXXT8wxKG5xyZWjrKxuDMsaqP1+Z6N
hOkeQi68QI+g2mradKM5LOB480otgqsm0NRo3BASCbX7wXfkSspmny1xSP0ZJI+j
iz+uXPUuTnjNj6+TI6QQxbGRTVptcTL8sWO1tKgdZCWcOYAEBTX016r90ft2ZLTi
8hLFP5kPRmN3z93hT4PLIvBd1YgJnzN4BCVEDxFeOgLruXLlzzFd149GuxFvjxtL
8MOGPReXaOjnrjqPMomp/v2zL94QqpbtPR5l34G9Bn96L0axCtgjab0hYtPGKzNk
im+KwrESqUQCcspgc6+qk929dS7qXz5a3cZ3yiY6/349WuKwKdK4ikwgJ1BwcALF
PgmTap3nSHGZeisAjv7AI/SyPwxQ2acUGGi2l+3TLaTBykOaUIeWt6U+DSXZSLpg
n09lAegcIvz58iJQ78ncUjMJ8reOPYTZ1gyPx1LgYnT2V8lITl+bmczyUKRcjN9y
98qGXV1wqxfKRK8Zo7vlZNlPulMpzMs3obYgMIJKUrVLV0ZAMlNCe1EzZ/ygIUZQ
bc1P8hdS176yYS4+Dxm00RMIPicdYVy513gGX22RVFg+bEuw98sHkroFv6AOP55D
8s/jhQcF+pjFApy3+y6pDAEFjvPqq89eIaXrAHWmmgdoRZyX89AXYA1DEKKnyGCG
bfUliayYWyfpm0OGwntS7f3kSSsTp/ppeJ9KPpzN95xo+sOdHxq8RjSFjziOuVN9
m11FvFmfHHeUVaUYYpHSq28a7ovOIxgfaGh3KMyG6QPuZcgSRGUz9awS0mpQmI3F
lY1m89xOtOC3/3pumuXD/zXbd3ySWQLEqHEeLo7PNwUUcCtcYuw4R+on/mj3cFSA
JO/89zbfKiUNrOnMXTtZ9hdhQe6R1dRLZ8pddukRcP1wLnKM7QfFYWd3jTI0Ylg+
sPtTz5Z655+pwinjSfcW7Kv8rH3xhVUIQZK2qge9ijzgeN6pxu+CgfUpIr/E9C5H
gW81FyhxlJ6IQdpzCiZAPyBebJJmjqGR/d2PiX06GPU8StozwpNqBE0aJz03TTZB
HxUNPOlGL3jM12xjqC3WmcV+RsoVKQcKeCuAJBpbDBa2ovCaLgeZV0odVZ+W1xP7
JW27A7c2BOYPwyB4MHyrZ2aDhH0ck86K8SCzObH1djzEeKX8XEV0JSSHXPomWdwN
BYNRoQtJkEJ4c3CBS80x34RK6FD750I5kc/osa39LTiMLT0OF0yDqnuCLXrpKsaY
vcNXS98e0x17B7mtN2AhnxcJMZXbCGXd6j8D9Hn5pbllg3Cwj+G39Y/uSrQ7/V41
mCXijc3XDYYvpU4QoEg13kYSql7+Zfajlon9zfkSc6DewK+Ad09ArnvzaiKjnGo6
ma5my+g7IzSlcsk2AVvnaQOoryGaTB7jS6aIHA1quv5eq6Na503RIyLlr9zF64Ij
4T3eVWWR2RIrxP08NhNA1Qo0elLAfenAFu7yjAXrPIR8jvMP/7eZ7tM/ZarRDS54
v2iNgPmU8ecbhbWSPvBxle0/Lyy0KPabfrJ++uwAoj6On8pbRGp2O5z0ujCMVfs6
uaUCqtxRF6Hf2Izdwln9IS/yplPoy2LFAePDTEurU9m+u7udP+kapSDO1pRU9GBV
0xLVyFBQb/UL27XOPPtKielbevY2AjiRqwGO49n++cxg6EjPzt+/MkmmiYHRtHIe
YURFB/02mLMbITb3IGl5tpIBdEBJS5ApYEZSo1G5FXcxXVGVLZmWDCZoxkb5Nyx3
c5NQaXHa/dicUOYGgGrirROD8nTew4/rX81XMrfoX7tArVuxInD+RQMIvd4GGpUk
hdke2o4Cht+RAYKytEBTLcH1xS3PknJKzqtyyXZ01I1ZCPdlwT6jYaO6eu6kg23W
G0egA1g3uU+xqqdlY/fXv2TjQPdpgIe9mTcl2bvWVg4jl7san2FZAwYU1yNW+Qll
LX8N58lyhucaFrL/EM9fXUOte62g5W+mBoU7rwd45HMbc1S80+/RQ4o+TRE4N6GK
/FdRvDiEEJrooTNThgkR0FUtkTGxw/7WjbKinQVhwFPkoKoFhLr4At04k5cSljZY
if19HFFbyGbOsM64o9pYif7P82XcWHY8erQ203OHzCOgPC/4Xu+UD8gTDifLhKaq
t1HHtgw+ADoyjvUI2enCrNyXXZYuj4X7EbTtuhfwM1vf5s2cOdwwAdg4isF6TlvD
pMthGvtRCemAHHv1GRVsLMQaR7Pn6JCfhWxj50Gmd87u2YvcfwHlojKc+FMaBr6n
LroS4zBnLGJlB8z6ZrptbhUzF0sEJpsw8Mxqg7HuZAL7lG+alFxm1EunzByP6I3k
/TyPi6pqMYfqVEDocEoGh3pYvd7QnCkETK+o6YWp6anVuyKn+vhGPJUuMJzodmKt
aujqjEIokHX6X/LoXeS9aOI+vNLb8wnJFrvGn4yiy0aslF7QwyQ+F7oFQeAxzCGw
L7Od9WtJaRAASj+NTlABJg9rNbi3eAvZYuLjEkNJtWMpEBMtuKiVc08/iI8mlQ89
iEMqxBWbkR6c87AZambuyqtcxWYOYsxqzk5PGFsgZEyDY/D0QjVCXYqhb80yPw7P
08S0H94z1Dt57b0KeD9I1FwmNMo6/rPCIXh62YVnMcMzQwwFao8V+d4PKgQCCRm4
IFynv+yKARzSQV/tenL/LJl4KPnwUfsf3DgxxBcvrtdtFTPdCvU+NNTXHltMxnif
0MEmSSvhkfJd5BhxOCgNqtRP/q+sZTMAKHH1LyM8poNxXnZ9KKk0uwluKciBTq9f
KrSYbnrnfPkak8ASvHMiAnwkTSmtC/1FSsNcw8YiSL70PoGdvC7AULi+bqW8tZWm
OhCjRUcW48z5CO2Wf5O692cr12K+hfPpidh2Q6lbgyVLMEnkmneccgtiwdFoFhK7
Xe4EUwbuN74ZI+2IaFH7LHWMERH1orC9ML8A5BZkRO6YZ0b+sjIqLGcQIaLBcAKH
KqZMtth+Z/cr00SOAuBut/59xOQ6swdGDgAmhqwHwIII815AQB3ZRf8QzI5UTEcY
PtuwkvP9ynMTKyOzyL310gJzq7rWIc3L+NsU03eB5rECdYfhLTpEKgYT4gS9Br9q
DsxwL6nyYKcBpi3fRBxc9nxOKCp8XKlIIfC/Z80mXUoajgxX9MJ4tIQq2MsY5s8+
k+3VpXJXsLSRPTFyuIQpwA4QQm5W74RV+OXdOMyf7qa8a9HmJlrBA+7kfVO0jb5f
MuHiNYnPnv33kpPwoKJQw9MYI63KFApF/I/EUWUg5WxaHBigjdb2g3g5+i63ZaJA
/cddlEsCBjaK9QaZsJNCvg3+CRd2EqBWAyPNWYA9cX0Y6ak+HPjnywXIoJv45Sh0
GWzDsOrSuwhdrjlNdo7bHAs6UsORuFnwQnTtrOXfB27TUAhH1AhNWgtQoEIXx+8d
4p9+AgfkwJSoPuFdJ4PFe4uQiQNCyl1XgWP/EzCUzWSQjPKfeO3KBhQJljec1JKL
uJjU3Cokm5AzHBYckOVASdRyKTnAWkt7CvgmlyNtmtBtEKFVTpL+OIdVRJNfp6yy
g7EKuvm8MS3f2c9mhoGe8VogD3La1fGJhBwlfaJqiyUeuzAgE/TxDMD7Urbf1Y4N
+vOUbwDGeyIHYZj3qu13vmn2xe7ouvglVvLUtC3gaSNHL97XFMOPS6cJkJcJ/0wM
pv4ZZ9ax3y9WEaWHlu54sW3ib9L9kNbZR4hbwUx9mhj9GHogoaelbELN8o0gIax6
deyqahss1+Ia311LnhVHyfXQHGfTkey2IWgap6DVWw9Y6kJFN9IAZWk3HM0Z21jj
e8TSNpbBU25xRhr/ji36FOAVwtu0e3fWsJaa8tewwcS3nNzDvQBIRVXeJOSvfH2o
GhwKwgoEzeirvY1n3n7PmR73h5esk+PFjfgHQawKyLI14R8loWUj6QC4lx+BhZf+
LyJDYBW6N+G/hAT3Sx70krIjqfzl6ols+NhgaZH8Tf+A+mTxul+oGwke97bondIM
JTZt24rzVGV+E86Vc01JroXg7v5A9kDwj3MwUcaKpVQDFuSvKAeXTHx6NsixnjYa
uS0l2zRZq+lixdwKyndRDdRRm0VUYY09o/Zrgww6LN2nJHGvl95RhBkTKmN4aSIL
8rFrhMwDTUg303g5YStQkrP9GVoeoZOxyCuD9nFaUz3SeK5Zga2NxqzWJyRjCFaU
q7lW8wkK+jJB6dk+9bAkT4828A1//3yFVHU3wArAbAmlhdYufFwneZuh7P9PkyJd
jWNKXZSW7HKV07+WQvQltQf6/E6DVGHd7r3wNHaC8KiY3eE0NaxuaXUMeF0+zPsX
p05MVE3XzojC4D8VvVI93atO0Snb4FpUA//2j9XQX4Iuy/tl9TAMv2kSsv8QlZUf
hID9wi8r5qAYb5X9QyJmzJkpsvjTZ8/d85i+g8hxrnrwN+95CCGA1/9KtYBoQ6sa
kT+s2pHvqyRwuwtX231UGOdZsbsRK805NYmy5FpZ9Jv2VmgZk67iADWmGrIN7EXs
hy4DQA/Mu3eYe7nR2PKtunfzbmJtSmzET6KSDbc2oXQq/A3+zWR/SiFEV6AKB4iJ
gWNUfQShBp4SqLxHy2xFwwaOekQLduV7Kpf4PNdb2mjP4EsnLlyiF5DUwkHX/1y+
8aen0Gb4xWJVi5MrQSvEhzhwAtP9PRb5WNFshpwQilLBRbcnY2p76s0bXVmZ3kSC
9/KDYB38i2QOvRow3xCiFrdMV6C56a32kZZqsQiHgVSaNp2jN7iez86fvj3n6Zbh
5gPseXCSoacuxT+1xg6KLo3nsTMUnILdiEYFvKcA7pUFS+l5sXcGBummH4VCQWZP
H4vL2gpHCfInO8Pop2pUDk6vgO9/gf685OzWdQCFl/bpotR2TU7lX4dl47wqhrps
hKUkIsSeqSxEsbdCH+sY1NB7tXI3qsgUFPmh5/sQzavukM4YD6ik83Svfnv3dBTq
8UXroYBoH7xZa7ZNf86axWzlkoGGy+Gg1l91CkBYV3+duvvmsxHosuKYKKcpvLwL
M/229L275YRFncidxEl5+nqvikJy0G4Dsst3ThMIdaQ6aET2yXAF/wuoYxf1qWeb
ttz5DQ2Eug9oa1+bp//C6cr4iJ2mncSs8d6apKuauUsONloeT4NZX0JwAw3A0G9h
HS7GDedHcd7mVRLiUjFFJdqwSFFUF7IwKag/DDBEYtktlcF0Aqacdcs4xV+Kk57Z
5I7eTTkTuIvQK15DuFMncYGyNUhisFu7fIN1T0DLYYmMyW0nhz/X8W0uCru6Q1D5
fwTHTYBkoCTSa2YYWAgUuAkufH72B9Ez50bpyNLiie8vK0RAMrMu4Dt6ACnbD+Er
ioLXiWM/zzlNxa+ZsDIzatS/PvOr5YWVtoAwzjyrpnjRoJ9N+XPz4ZXhPNjhkZnb
oZaQC+1/kpMTbN6y3XKSsfOpBkYDeBpcYuY65QEq2pNBvNF1dHdI4VQ038Nx3ISu
SMwqJQTiA4cGW5pZ+AdpHc4DK/hR4BHKdfEs90tm1zJgEcC0lf4UIzzYioVlvSfs
nDjmXtC5MsMKuLCR+3O1qAnBk+P/hhsIq3kR+Jav2fgFOBtvYZfVnq2aHgH6m947
K2WgVww7qk674TJo9Z355ncD8WXY9UZdmA7pPo1BiDc2r0kTHKs+BVdghEuBQ6hg
IqB/H7kBCjwHyaXWZSi8pJmPLRUSOXgZv2V4qXZFBqdd0E44OhHtFXAYoZFIrZ+J
Qg353tz/zCbWApGFY/+Et4Mkg0QqZdRZpjwF+dOdKshfwTEmrVBr1iArXUe/tYy8
Rb6UUKUrPDcl4NEdPhOkBXGO5Byc0lqEBgQxhE/XBl0S4JxJB9yqOeHzeL6Tntlh
yffJCxLGvymgxT0SbWOdgZ0C0VfrlOTkjlEeGU13tzvSjXiaArRe/vXHqmPvh6jX
G41IyWQQSHMrlDQOCnkmJw0WEhpqeBI7uZUphtKIly9QJkoDTIQWTtzLfDNJlTih
bIHypVoM4G2hYPYV8nUA7ptM6QzFdNnzl7RSfA7MTdhFpsGvs7efQLZ3iaRa7KxF
gqZ9yVsFrklZgqcFgeQMcvk+Cuc4Ke53Z+8QRHFzR7W7/q4BefSSyJZaRtQh6JFO
iRMaoEhbSZJ7q6d4EDK+lUmte9YRqHEfNnJcGvL/rzY/8pCLxDPEHwwUu5c05mtp
49zdeDIeDyoP49j1XPDWgb8KnCTGWA2gWbSXiJxfbMGLzCVlyn2BWezQXEFbKdkp
BaxOjhhEnjp4bEPWNZwYRZJwfo69nwHiCmOEBD3QePs80i+zcExLLRatAB2GpJ43
ffFhO0DBKWpCnjbMsN3C20cMNJtA6JZq+ix/yYaovBEsIZmbPLbzjHJIrOSyViET
omDUd2BVPWP4hGHmroF0Xl6sH5PZnUVwEsTxFbeI+psHGqHndN57rabcCZhDY4JH
9DyVttWyTDTAa6zKqxjDZOGlqv0iNySpRdaNhVeZtXq8rotPLlEhgLPmwExCmY9F
1ILBKPWR0HOcezlQMjA10P51E8amLosdvRDGU8e4JEQJ4ISFXtjgjnUrAm7Tvf8J
sBgXVKGRI02/BS8gZyz02Uv+lVa5cBPFpuA08ynfOxLhzZZsbra8F+xfSN0ljaCB
CeIMjge+AHtvjDDKZH+HuKtjQQgm4oVlufttV8QqCbV7dnkEqLcfdpCSgeh6j22a
cB8HdqriwstGvrcGNAziG6/+Z+VRbcfmDcXueUAXxhxhA7DPB1xrL7323/rKtBb+
JW3eANnuKrtZPdI+kZP1JOAiDzTJJaeDM0I0he2NhCkumBwE5eVToC4pUDX6OIZ+
8HNCho4PDzqzZd9M9AXW30C/F3hV/XfcLtwGUsaRN6TCyMx0KN4OzU2IEotmEBWu
qnkcZA1XfuY23bcXY32PLJMJRbpfWbFLcNApxbz1Wum2ugCFlrsRinBoYuIJrD13
vcZLIOFdZRIWmmp5uRBlPXW+R86y+gmOwGFYVT6OdS2Nt6goqhM7obvF+Mge/e29
jwVKgYSmsrS8aB95J5YCV1sGJEbLyfIPBVkzLD7BdN4pHlV8OU97nAaNcxTQEs9D
4U1ZartxF6bb8G2FgTTHWjj4TZjW3O+k4jKIAzqOFHMXUZSnLWvAij20A7T++VfU
100Ulj/jx/+Cb14GB63B4NXHwn/HKlHJB8aFqgAUIT1qxnOV6gi7hsIlKViePWd/
6nx3wPDTcIv5ifmfctW0ctsQZuBuPDoQhDOZaHFsvItJr7uafuOF9bQFeD84Teqq
4k8GXzG6x2lD5uKRRmY617G7djZaeUHGDC8KMUWJIGPmSnZ/L7J1X9gQn1XQu23r
zI/Yx7d5cmSwMhgDXMdWGi6OcLa5KDBIUXCpV+sN/B/GElIehl/llroZ+J/948qd
Uyg2y3LaH5Vt+TefD/aOcN43zHZ7/S3JpkuFRTAt4nv1dwW/TRN6JpAku8VqbNUh
MaoCG3PzTQ+HXYB6sdk95owYEu91wIzzudix8kgFZL1hStPWtbWgyy9B9RVkI/z8
MjzUSQRhqzavKVD6efOCS8UJ5HyrPCRXRpl2j2kpPGx2N6IOLESpmPvH3WiscjlQ
zn1p+KkhBMjhHCkYUwdpTHmrt6kCylMpayxT40TFCbKFLmQCqblZvFawRxSYTC9U
AyHFJ6J6LhiUz/KxIpBox4UmicobrlV/6DImFuy1bwJSKdt+fCjptGSX2h+lyeAI
0dFsu6jCgoZ4Jaa7JuA5hN8up52Z/9t8zIf80tS0Z4EOnk8e2p3dcmsAuLiZyTAp
HoU9vIR7AfXG6QEYQ4PlksypNl0jknQVuKlVcfKPQoqraLYiBsUq147zYciU5Drm
ZhakIVhDQF52xhpGBzdo8NmpXXrM8KheStoWEmMIJhoPIoUtNkYe2sJEUxcAvCtk
3aZW8S5rJRp42pLVNkLtUPdJQ54FMFQWyCZ10DmtXLRQXkgDvZCW77hk3TRulj2f
/UpbYknVsiXMjWrUkrxMamnkCv9sT1kyytuacIQ6uvjPtAYfvTXLMdW47TvWWF3e
c8mnunJMaXHlVtH89EKoGM79/NMeeV9anNQ40O+OjOX/4EV7YU1uY8s1BXHAgKgd
czZqrxOnYeSjqmD4ZuMlcjptS2INNK6u3TFebix1DqMDQweRuNgEdexR40MbRO59
mY/V7S85cR8Im7Bhs9jCGdzjXOgpj5JyhNlDyhSKykbzMN3urPMfwu2b4dazJDb0
rWkQYBvcOyWS6QSBCMaf5svQ5WHTjN90FGvTqscz10QCWVjG9QLnZ5DKVFra0tuo
t0REX7DDQwkjh9sCzBeiwWWoMYz1CUrqZxcyFu62rkHmcBPI3VGyBgFxHySt6VmO
yo798ek01jl9h8Dia+EFTeXjVeIc4A89mtXr2U1W83PoUaHpKbahdLqkb+J6hRIm
UKnX8ZWyYfhOvtgt7TG4MaAOET8jhg8+jR3+4CaS+Bv4xsW2F2brj3ZHN+/ZccqL
iAbHl67afLRMS5sAEY2bV2Ruv99e6oiB9sXSWsleSe7QxlDORnvQXme9OW6uOvF9
ladKJS7QSfnUX0F0Crl7XFS3/lNHtNF7VBHUzdxOuKx7wkWRq8Xup1O0UjOQM3QH
PcijbUQpbPbIanDdDoJGDozPkiVP374lFZTUdjlBJgGZre4xnLwF+da3Tfh7IAgw
AhI+NRkCN6zG/SwbjSmawezPPsWteR6A+ENSFWXSBUuUFYgblF4qPau0F38Z+BuH
sysBZmPwdqrPlz/XHW5joC4rI1g9czM/FYU8CpnJ538V+YSZXiH6/KFXA2mynYG3
T9rjqh6ZUz2bnvMq+rdzs/8M28XNT6Dnp31zNM5MeZTiCV8w9c+1eYWU/4aGk9en
HsROHv5fC89bYK9P01wALwqzi339YtPbu3KsXqfVYBexRkdBLfBKouvnOUzdRYgP
iUC2wYvVs2nzWhTICtZQK6S8oBBNJZm1+1d1CaV9DA009k5c9+2jY/xpw+IthY6i
zTLvxYIzILRsPt0/tJkMKrvuLjoDHNa2lcJLk0Eb+JI0JXerhqp4SkJ/gY0wBew/
LH2nRuiMUb3f4Delt6jf6nNhxeCLvOqSsohvofDKxsLqNv2liQGV8iKhM0aj0laR
t/HHiUj6TI7w7jZWHquNuwVwT8wZG1Xj9aZ6O2jxU1dqFcNuCU0U1lnE45uaeV2H
3ht0oh8NeD9F9dDXiI3saEhLnTzQcv5OaXY7UFmKq+stIE93e3oQD/rXNQyuaV2y
Z6d6PtryXtaUN8njhqRJBjrYXetr7TMxtQOWcYyzgvkOZW6CytkPsRrCvPkWYO5C
VJP4Trx7hUg2Awjb+uqCWIWdLjAWWnCioorHhV/x9m5rIYHHRU+iGzUf9efS9A5T
tMNc0heBt6WsaK/cICNTLhZR7HFk/brHMktLNBMu6GOJbPSgYaDrZYsF6YRYaSZy
zN+F9LIHWRM0ozeW6Mx7+T/IyV2CcALWAAOHRiG3t7kZz/eqLnWWmm1+MnhOG0YE
j5jGGwL6OfNhE15bKbJI5sr4ZwP4fnsTwPQkepbA9kvluJuKgwyRwTwSPTgVPEZn
GhHfDEGE8sFCx0FqVfb8Uz6v6MxCoQmlmDc/eWkWKjGYgUnz33ehbZKv2O3q08dV
ED6qZT60/XmDp5ri992F0vCEcKLfLls24RejNjyXvoD7zNyfjUajAamsinmXCpXT
9GDkr1QKwUB9LlUDJhgbHUijjNpH/iR1uZgWsTSJOn/rcABAodwJf62iK1+yXjRQ
eDCYPHYLtmYIt4eVfzRScZ0cW3rwa1jafD8tRRrCjl+bj3J5OE0l82SzetIOYbwP
OlXdoEAp780jGnLiBNFF63XzhaKsq/1tC76T5GEUR/YcWmuUSiJZZu3P4On4gHlk
rFg2fG1pCLaVV2lePirSi1kJtooiLHR6joutXrsAv1errIYEQ+cUG0ryisSCD+9t
aaFNXw7naHUmmYA66jAXxYvJw7E64Q0PvPMfXbFMguyLRK9sx7NGqjuloaKuMqEm
/y8FZYwmWL26wI3D90owdDBWGo78/6Cp81vfUxmC937/nz8/iKoZxyeZfM4X/BCP
doC27q8veiM0lttV0TE+G8yqD3oMv+4H6nZFM+cKOPV5f671vDfJaF1fphed/93V
QoQ7fSjCbNazV23cA0KJQaSuLtUl67yir12lASVX6KeapY8RmtLSbMSB7IHufjBg
TZfdB8RIhpgst8i4aXHAXjvh4kWNbDDHsesaes76VQmSk+i6yOACcx5qY0BfFqMu
HeVgaCw2r9iOzbDMdAilU4rDTpGAtKQ96rLe3VTvqYGufigj4bgMoJoB8KRaaVq9
7HA7U18pfp+TEaL4A2eBAMLvJd/h9MdUJbgeYBUKLBUDZvQa0JKa9jsiQ3B7Zh71
7I0Mzvb3g1EPzkJInirtthL67NIYwAzrLeTPFORryZXdAVwOT1utSt+Yy7fREEfW
/FTGde2yuLVAcEI6swoFB7+4poJFP4hK1YfjM6ora5yPMsfWpr8U1ZiTD2moJVGg
EU2LSO0YwKPUfN194eRThhd3H6rQK2j+1pvss4mmRrvzTJ+J9MnoTUXR7kJJ9a3k
6ph88GzjqVBbhncgjLi86Z6KPMMbPaF+A1WDVpNdc6G6uDs+5XHJf/EMfpCiqrfC
6/uBEXtiC6WEUT1wN98uZVe3ROGnPMf+JxQM4d0UwWsMfdxdCFwcf8LrPVPZwEW1
EeOkCP0nbpoXvI0CK77gd+XKpGKqEl3NNC4cUJZ/6EZTh5t1FpaTcJ2zw41iLtep
WA/i9gBNSl/25euUKM0dYEZt5860J3rBvj0A4+XkPVcxUgR05fAYui9QNCf9m+PN
xeKdYDvMdthKzMtO7h8YKlD6XTTpxvDJHiTD1TkMqRINzPuB7dJT5hmhFmtLLOKg
LxMPlS48UI42FAQBSNwWjG7zPzUm6g4ZQftttFRaC6UpesCSRst34TCv+pKeaHda
8nMtaoj5bvs0g+Vvzgh07zOOcP+ZxDdHcJOYd4JPgpgHP2Ze0AyCWj+kgiZqhBuf
NpP9itgemfm3NOm+S06yS/9S1Qf8M3r1aQ8nzsg3wTHfOzi/aiQsfgVrL45I0aE4
PdLifS1GJDFlWyPcS0x0ceNkRjeGjPgNfTWonNnPUyqIow3F7fvucIP0evVA0v5s
7IilWEcD2gupPwq4xbKv3b8Ga24KbQBGh3xOjKma/3xD6Kfszh8mX+dM2j37w8P6
mFtkfVRoouLxBrpXAggRZnjzCWMuhn14npDHI1Vs2yM5ENjoNJ0PHNnWIGCrGQ92
QKQF7za766j8fusobNyJ+0XJSmqnfeM7yUcOZtFju0/4uByO2avjE3qgXKFmVwYV
+Ku/rdafDRqQK53pnpMdBBIXjPQno2fc3AjUMkZ7pqIAJedMUq2GMrHDyVKxZwEh
oLaC9VimsGyL0FUrXt+wasR8FloEfUZVxrBEWUvD8g+ersACB74rZvPejMZQs/nM
a3vY6W1zAmUnQ6e1rB2lkrDgFjWn9/ebiPqbsTXbvwbS4vxHgq65jS/8io3zA6SV
CYw2ZpeH8mkBGG6nk+bW20VKZKzvP4Oln7rX8oLIC4z8NIJwHEwiS/QZjnTFaK2V
IwLX3A0D4/WA5u2LjY0xjxkya+F4lKFDE7fU7MzgRqT6w+IQLlkwO1mocsn0hSwM
onK2fUBzCAxnxBhCWz2b4d5nWYMdDZR6WPFhDp/0ygUoThAuaKnjHLgF3Z1ZipHf
sU7jHoNY/E1KWzWIsUNgUvLnhhQ6QlWYtV3XnePOtxeuZY6SBctzPQWZrjsgyeRt
tRTYTFBu4RBk9AXXXUfLUvlEcqHcmKWhLUi64u7291FYMZLBzJL8qSYjEyYj/C60
xkL5qjbgYqWfsPv/WzCPhl6WekLTBUUpgwdSNadeKqtjAlKy9SQEtDw5PfyUFEOk
/+QfdGnyvuaF6nzn8J0TC62JZM969fPAfoUcAnzMmOHhiPniDG68VKuUx35c5GOK
EOjccUBdIUgyAVpklg4FD0atlZwrMrYAJnKIFJTYlqTNre1Ykcao880yrvWkYH3j
p+f1oAppXtwcLnV8J/NE6W/MxrQel3GGOEleo+xz2BQ/ytZJoMCQGJ2iRaKMTD4I
d0yVPczfRwQrtwzPUnXKCpHtWngID5qfmKkZx1n3s+QzNqcCguCjTcuCxPbXJvvq
HWM6B9E+pPCOCfeneELoN5lvHTNWpxbP/DX6JgHv6Wl2QFRxisgqXioRs8LnRVkq
Bh3ZK8jTmcYDf1cdgnad2E6GK0jmzJZyBRTc/NnKWYlzXJvWfJd5T6FwBOcpHxKz
WnzranjCA7REepPwNF4gvTVOpARUHIJvnHujnewTrjVFErVWAnBXG8muW6Dj7swL
4IOzV7YEWG0C1Ueqo9gMCFjpxVEt4yVdgWQRsFcHlJKCfQl4Bnv4ApUUFHgDErXd
P+qxWakpBSz4a+yfsqhcOecKIjQcX+CYrJVQX2mJGBK0mBxV6pjDoDpb2rGsDy7C
QmUNXpFvOwI3YWE5xT2EduZJYwge8r/M+UtjfDE+tl/oMMFInXoHjiAsZejvkIyk
ADpI4pt36WfUv5kkTQId03wvfKYmCGzStE+NatSIz+0EVjVkOU91IoJoZA0JrOw7
T2EEs0i9ZZnXD5qMzynInWzKx4/p5ABOLZsi/7JksXFf9ucznl5HrRivVIiQHXD7
yp7ml4YZ/N4Zs1AeYs59KuZRwQjJkArGJBvPvVNZTQsgOSuf+vGXiX6PXJBNL8un
XZ3RGgw88SOWtaJvYDDkQCXmb+PKNZaMMBdodaN1XNextSwT5vWCMMuVkxlCT2Jf
/HNImZjX1MlMpSW9PoCX17lxYarrgsQL6piY1c1IbGG3YJoGAWJboqbk9Z3tEgbu
x+mrmC7+kqumZd2enVoTYNP0CXDijTvfpDaIz02UA7QpEiFx8aNNFZjTRAcdi3iQ
mpDBhFKr+4jEPbC00+p14iQEQJvzEkbu5iiXY1b3UUntStykW4nEqQeMdEdbqbC7
XwUdxTEqjWvYXAV8gdun2i2NUIjoH39LBdWWmEHhN8rI8FGILLhU0lAMeHXvlh7g
LGpJQgwArS1ndTOtAnwQBoP0uRvmPjpGRxIoZHepbspl9dd3Eq9RCfl58Vc9mCaT
qFb/c2epJ52wHjuZCOo3i49w4CLc4w6FsCGjqAD9KHciN+wQL0TI27V+aDAqi/7z
dYUceeoV8GxVGrHGuuuOnqxte1jrPtJDp/Ykszhnyn4cd5aIdJNvEYNCrkEEXyJU
cWCbgJB8kXVNCNHLJ4jJVDz1il0U7+x6yAAJdJm92gX87yyI+8KEPWl066kbSSNx
scqMO7A1YlA9fTRlkba6IZayHace0Rs59pkxYibrrqMTCR/M4lA0HwfDjQFD1cnF
tus9FUT8tya54/tGApM/04yqMJ4i0W8boA/gDWgf1e28r9h8kNJalg/9+Yn17kJE
dD340zYY3vGidQ+q5MNe1dKmiKiFkjcJAIE+587aU6UXYmYtKK389gIJoYBqwuWH
f+3JfPvEY/UZiQKf7sWEV6tla4rX1AJUfJ/TxZO8h1pzU5IoS50jkflvw79s4Q0N
zu9ZMRGjMGKn2eUijc0bHdP0d3oYuKn9LsN/Wcvl6+5p9U2OZegjBylJsmPTMoaB
euBf4T3PU3vVvrFaxNGyuO0bMT210kMIWZTlBreoCDTv0TjVB/d/kFeMLpDkVHVP
KS4jQYo9kPLQwbWHKjguTNrwy4DiMzcEPKXCfI8rWdQxS+okGEHVl3RDd9qm6FY3
+ERtfvXEitYyZXKExh2xodAUsKOu5jmHRQ2k8G9TuPiyVwJTu19fPHqbftQTDvSO
Auk1VcoEfIB0Hu6SfNZRiTAlLU1sSR0dIkSmt7ib6T8q8DjwfNqO1AkprpD7c4z6
EwVaQYWzcJrgvONAhaYoUSRl0CNdfDc6047o2SS/fnEHwMXPRD6wQgxjaPWpAIvA
KtgVMSoJ7oNGpy3eeo29T+AqdFXot81WDrHLOvyzk2Qj46U062vZymrNR3m6DBot
DYMZeiBSLhhA/XBmQsQzdY23bog3lElJJfVC8wcfvfFkem1H7Cf7tbuLln73SSV2
b0T5NZm4W+XHKu0qFSsx9BzBHXD1eDEFVwW2Qz1z+HOEVXMSMVIrLxNrXR1Vab56
ZbhzCGXopCE4WmLlgLcU/8Dr0SQ9ZyW8/FoO7MaYsGwh72k/dUltFNbHWqpfQxnX
joVOvsK0PoGHJealCQRiMI0PRjDDatEKWbcNQqidJ/lPLTu4HssLPmBQjdZoWB6o
ohyWgyouj0tvbgybveSJiGCQBVKNHKFyqCW7I6QURs+q2ALki603dOxbPaqFy4bM
TKXO4ODI42l3SIbTuqwki1qNFDP+H/uolp5aL1zepHP41EVfbnDyF+tqwlbhwHFd
3VdsOLKh/T2H/7kSYDQyQSNgP0MSLkh/Mz00/LDzufd0JEMuUil9+oLN5fzr5FL6
J4lrt4ftsOVdPnWmheJFgk2sjA1BDR7GJpYUQBk7f0j+RKsYqvM1spcdAd8D6yPk
EhtWcRWbjfIM4zmLt637J4JSRC7c8j9tXP1m7HoMBVNdIadWe5De7hLQpov4UsZn
LgMWlq61s9EpoyiaNo3taT0OkOEMFVIHOdeFOktHP+SF5XKSG5vOOwZdLcxXhU/Y
mKGNyZf4U/Y4TL+KLQn3yFLTXFlO7O/YZqCuDDUpJWhHtxW92QSsPTE6EzB8N7hC
H8X0KVERvSOvuYnbrwxxa/KxyeflpkFGStkAaqQy4px+k1v1pPaNLMPdbj7WP/Wq
L4YgEAhNDVw2NDoPzUnaB7J+5aiYiiwntpg2zdjMrEZ3c0V3bgwLFQOoOho1hO70
0WX+iz2JQvUaWuZjilY10supGxf12oMc7DgDi71OYhzwrAD3utEILLjo2wEARyV/
v79ZuRzr9vP7/W4PsI/9dy3FUd6fcsTPIRwgR49xQCLkr+wgYjBo2mZd/IMq6rGT
IF+KZGRu3e31Ooz7XOy+AXb7UW1Jc6bQI70m1eBbJIe3P5Zr3ckXfJBrXp+KR0fM
qO8ysxtr6jM2RoQlJEZ9mZZPcr3OZl9nh6Qk1q+vM/RhK5gKTME0y7u3v0xxY8me
nACtJO0UjiClLGY14Tn+DkhZecH4m8sHdaA+/+oZcGcmtxvXHmfkXzFmJeDKXE2k
y7khq+7cC7aVKZmok4QIdx7QVgRJl9jvR4Qgq5A9F/nF00PQ5FHZRaZfU2x6B1oT
oALTWsNCPAzm37ZzjyGsweV7x4QTSrHwM8EdkcpiMf4HaSOWTpl2BGE9o7WdLE9k
TEZB+HcbjwakH2R5ve5Jp8tZefcORZ7U673pfoVk9H3ozeBgT1uTUFRcpIbYmEit
UFOnvsibiRGUqzDf8+ULIWn6MGuHXqGro+Sglt/wodsNvVNUnN3L8IO9Vh9c4Fse
53XqCZkXMNvYaPOyJuV9WSS/jVJ3g2zRX+WdHuDNJS36AG2EIryt2cbtF7/PbPFE
Ls1PBLb7VJjRjx/lJTVUgH/Ql+uMIw/Zcrm4+p26viRW7EHFRjc2ut+z/oWZ40yl
GEr+8Rg0lkkk5erOl9dLEg78MfTzH6YTuXicAs2KcDGcn0aK5hCYoSOQ63YQLQ0S
5Zgm+x5ovs9opWbJJq6DXV0zOA6bqVEtKRlTNhxRZYOvbU39ffiZVxSMAs6KRnqQ
5xIU66YS91qubjNMzlLges1JTKEXmubcJnroouQtgfZ2Edq01DqEgdZ3a0pfihTm
U9FGrbPNM6wmeWqrwYJlh0bzl4B24S86S/J+xbFdSj/18xlVmzCKtx7nn0JqMC6Z
MMtaLfbCv1NynMoP8EQ2h3fSyOgzgupgymwmkRJMIp42H/zwbnocx5ZaRqms+pak
kS7ONwDTiqVlsZ15xiNACVeL3GBji2TG5Pwf1hSDWpB3DjkrD3KJOCDW6tMTJPEi
66VNSxHG6FotgzgN5aCf3ejLBsMOT3Cgs+3JBJtvpcIUJC1nsDGQy7DQfVodWxz9
+sgnfvqy4RUl9yQ2zqMUyJg8rKIAQEBZ3B53vlP/7FwjTHrGprTxr+A6I9P0BGIx
zIOm9oe2zl3r7mA7GsHrPpXAYWjAR0TS7TyrzzWd/mRKDKcpsxpp+axWgNrXBlv7
2GrOlCk/HFk2/ieSNmtsoL2ayPS+6BbMw9IGzK18Eirh2Tf6MB+nrqL8k/eocR/e
UkOiYpzJS9TKjfQvCQb5EQjrtV/4br5ih7vO3191zWOuxnUCtQolNVWsgYGQmTI2
SOQXcEGqZI7XHUfWGs32GLgX1BAL417Wm8PQ7fyyid0e1nMkAWBlkTneu1EsguKC
TJEDWXCYHrHFyssEFvanNnKNp4J6vaRg8QDgZ4vrNucohJ7Zb/glRie+yOrAjz34
I5RCOGD7ITTpdvi6OZngXHIWbGzAp8d4dO17GhLqIbiDMFr9U2oQsz0lwX8ddSHm
qWdfkO8KzmCdxUYdTHVrj+H4404dNL3eufPcljj5mUFikPxURC3CIeCj/JyKSZlt
K8QhwaCCjdippH63gVMGcHEh6xQEPNLOkcTPDEGIU8WLX3d1GfmepRb+0dqHnLp/
gJXbABUUgcW7joElU+0udbRoToIQddgBeLYyeJ4zuN+aP6j4m7weGxpLlyVG2pNw
rH2fNT0CpVoMWu5bX1FI8+WoRlwJRJshgW1Bq/WKIs6WOFNe+zTW7Sj7XwrGG+d1
bP/U+ILbg491Eb42pNeUAOm52h8zoKMEBEWo9y1aaaL/Y9TNWptAjm70FmGHRE4c
U3Jx4b2T09740BaBGyg6UuBEwnQXkVWkADnn1yDhTV3LxtY33Ov6MJYlv/MOJ/zR
SJFIwSyO/2mhBgMC043y29AD1dX9S+koU82V8cEKh63XWRYYGHIW6Q3hszSmiskc
orLcU5wIUbs/qC5ygjE4lR34SxwZ8yconcYLPvOzKpo3XC4SdDivgpkZBh3XfVCc
EB4Z8qT4vKpR3tQkfTU4IiohbVMDkxVmFmJS+dANVBg8qBxdg0PgLsTrM3jq0G61
CeyEsROLAqG410tkyAd29k6EtClEysfgxsXlJ2rBzwx7tIzFpC/yeX7/uHxKyljg
Kk4rfvfOOzjNzuj69quMn5XFxfVweZXh6CgFmvVFep7CYwjfarGLkBCpH3TM5/Lj
XYKWY2H9tVoyhHK5A3xyXDM4E2HKaLEAHoYzVVvtbm68aO4IQKiP9GsXgVnnvm2m
4bVme8SwYZibseNxLxThEBt/WNuIxhsCm5h6cqFUvmDomATO/Wx/uhLw0Ns16OzY
jDdZlWClviuWUKk7JEE4tyOHVedooHaJSCMxhThtrjhrRes1V+xSK8UOyIZxVhB6
y8Wa5UDulbIbL/iCSnBpWZAtb2uYmn0Ic9IQYWpwNJHZvQmrmTCt7eImNjGVcz+f
hy9GR8mvI6V774szwtXR6DeL9g/BS96d2IFwIlC7MBY8Nc4X+BB7YXkRGtxpj3Sn
mgQSzaqJU3yEo6jn3tnpjAsTLgVNWXPuehrijsijtjIQAcICTdMGmjmMddWGI8CA
ymw8a/WxCLrLrKfgk3KjFQ7IigF6nLuYsj/Uj/db66JcS1cyHy+gOprrSu6Woe6s
K32ZpjXiKFjQmFB0d4nu0i5t5Jr8VeJNqQL4bVUWZRQzA2Sl9QzqvULvKtCOh7wO
AZYrpqKs0gsiPh0qS5fUnYagsuiVp4XBtzWZ3vJOYB1Jcwr17eh3tF7IdSZlcoLP
060ay53F1A7i2C7UNIM93BvG+oIvE2ypNAmgWsvJPvKmiOBhnIvWqHUlgLNEhVUU
h7bsFmIHqsTMSGS0vyzxSBuuHhOnFntv5CCQkP6OO95cK7uiHUN7SZjA6Mv3aYKI
JxJWkEYG+VmoDR903MJfwBAaNhJRCmxPLrkYquoym95hmBsxqSVlWOr/KurXDaWU
8w+1vgNWBGjMJ9ggoM6F5Udj3qIfFx9IYzusNHYKE5n8npm2MxtY2/YHzwOWxlc/
CXZVVN165Gp9e1vS6nrD22mMkoKzJLq9/jY3L5CJwtqkLS7BFAEHqeZx7ton+Jm+
YFMMbKA1Z/Mf3r2iu4hDFSK2XnvkOtrr9TePzsvlhaXUmvfAujHJZtqOUEgplFDq
sxRKmUVWyfStd8IsRtgSKrHWgFgHugWXd1Rg4zHbL59c7qB1DLTqmC966yEoS4lW
16Twnbmmr+TNsFWMsews41xe1wiQ2lVeB/+hwuiBBOK9jhToUkNP2LGt+CLiQWS+
hyRRfCJ/5XfRgItnkhYBjIfdHFm0PTIoclkKMDZqA+N1Ycl0QWUjEhaon1qlk1gR
pon7GdrJ9KKqFu9J0X7itQS/vnLi9vyCIh7TF73cIixsqDImgpiFVPUK7ceNAASR
Ps6OaTJBVVTUuVIoemBQ44npk/AUCtW7PO3mWA/S0yKbk3i10meUe/lY5LwwaygH
yWD0+KXuoVgcUu7EeSIBDb+TpTc/wlBUa8fIq2tYtw4K8RMdVlR51GfP9rI5/Vbt
JS3TLVfXGiU/AGQOGW36BM4iS+oBJoK7qJeRxLiLRvucjpsTkCjZtYm9buuU1p5D
9clqeTVwtxtbVqxbwgi7DUsD+k/374I4xeXAD8GCWWnmXufRCPG3vLdtRhPkBNPt
pmqlkYozWYEjTd+kUrz5MfD5AJQQEgsi6sq8gli7SAPeEROxOj2FMTVk41K5wjHi
oxDN9SMVyLWSzhgNZKbmthiy1QGiFZLNG92RQXRQHCTLfUcXO3K1eugkHJ7Gmgb0
emjWoUktS7UIuMVfO+hi+vyAV+PRDpGoiFWFFUQ8j0if2mXta2Tws0GBrXrF0JZB
z104f+7Jffwx+PLTUlO5flOCWO2T2mrg2RTeT2qux3JYN6EKQ2xGkP0gh41UQU6R
zKaMt5vCMKC9tDxnzjc5lV/NPr2XBXwCvd/aUqlPofqZR/+tmMOWW4sVN9Ekn/nX
OCyTfdEn7N5qNqhhgukKcQvsIac1ZEBrUOFx227+gOt9H1cVVghhFhj8TTKKc/oL
Wqi1ev1Oao9HDYvrJKu4kbl+XY5aLtaU3XdQYmTAH25Qhy7E46poH8sEDT/umfPc
7BxjV4bR/++VZAMd/uFudI+w1XavpfQC2w2Gsrky8bE2d7syvF9ZDlAHhCxq1vVp
1aDQVYEq1zTYfHNiGaQX1jNq44PLE/yztQfQ6ee/l65bY1XLYbNp6sto75GgOYCy
BUL9UDs6FhfJiBIRk1T+GIXRcokC7MpO7d23kv5zhp/K7YsbkstxDYStxBoLk8Y7
H2h+eA6z8rgWkgI8e/BsvuvQGcy9eTOMYfK40GgDdSNaetmKwaEU0Yi0SwcW1Oqm
amGnrdhtUniFkDjbI0Hge588APpArk6QGXjEeEmefM7njMx/n7MBJIEWNBXoPWoB
vTL5jCtWHcCSfF9udkGwnux63/oYZ6ZIyJkMuFfcazhm3y7jrfLe8mFvbudU/Wfh
j3uDGroDzBd0KIr9KaG0fr3uOjsvjYVo/VuXQadP3Myq2fYeVtMmOkX1DbOm/m60
/gcnpmalvZcdPSQjjPhfhQYSUxXxhjIM5DFsjM+ITl8G/JDcQcDMvqbTqXYRr48s
rBAp8Hrhvx92ALqS4ptbPd2pavoxIwn/yLiyBULs/5nMtni6hBC0eEmrpMM1+lct
Kt5TVZFg7i/4o5Hfm73BCoc4YAQT7OehCILmPjqUj2B1TCMg8NSTCF6cz97hV5ul
Zkxc4ziOMImGIEMm/ZInu0Jv8Ljt0pkCMxWQ5v8iBnQMI4B5CXIHip1Qf3mGPTNJ
e2iBKiFIWAJDUrBW5WcSO0HC3QRsHazuteNvc0JulUqdhP1hLiZobG5tEU3pY4Da
tHT0IduUguvVuS37wWdbywSodgp6GcThNB3qHUR5oUfmb14g9qP7sCvfTxyWO1q3
71x8WsQinteCKsOOvFpq3pdweKK7FB8bDJ8/XmPK1Tn42D+9tAS89VdFa3n4gipx
/6LSJTyf2RYh2wX5NuQJ4bE9f8Bu1KNNIrCOhd3JrEf/GtMJ0LCNJLnW+EPCJasD
I9+V+iNPqEuhJaKSDTPqXVbtOmZ+LBArAw+Y/oidgg7ite3o+7pUreKsguQ/E3HF
jxVZ0X7tqsQa+Hv4T4ut710CXIEqV0R78IP/Suw42RNXHvROPY4xozFjS8+8Vxhs
3uPfh0zVs3pC4vdyqxPqKiqv6Sn8qNVHDOUnjVmnX9hzTSIMkF1oyN+mC4JL2jiL
rixmZ+wtv1pccLqdo0hI4MLN2Ee+Gnj9tj30VTjsBKC+vJBFmBKFOvOcyMswlJgJ
yVPus84tursW+mtGQyPHc1WiL7tDvCfNrWfzz+Y+7fINZ6UupPwdHbwnnsRnsrOs
oCdPbhvLgBh95Tzzk4fKmdXOwz0UXYoGVELSIfEWlteoStsbMrJbVFmrGnyup1So
+dWUX3rfncd+a5mE0cAsSJrC7YVH2AZos20wnMgkuxNnqMW62ivj4ovruvRp+gMh
qWOh9RQnPAsSfnEgI6WH4vFvfkmV1Y34olbn0DE7KTo9SVuu3evqYWTB/MqmHYnA
anS/QLPjypnOgBjx6PrfB0Jamt1fBQS2xZcYAdPj0l5AVYBmtOUsaexVP6I/KMUd
O2cGjqIeSDRBQJwhTtHxBjcrmwX/7ASMWaf+4+5ABgq4fhSl4rPOEMrlffip95F4
ZBqhazOAissnLh4qzV+UTMn2j3Jwg8uPpUuhHB5wrFAbKRny9uGrGt76SP7kZp52
IECzR5Dz9uZ8Jo5xlhfWjZrVgm3aYepKPflFpUQPxkdx0ZErDjHonKVRqoBZf4K8
D8e7VWQs4Ji0n34FktqRoboK2mtwtA9vA/Qp52UPkzQClUcoeSyWkhX8lWZYHyCc
3aeRhxoVNr8UQLLslRF/YxEoPXhMjBiKideAErfGZYKZz/VAjMjn56Z4eXuaWup8
0nepUHt6JvNjtYfy2lHruTPaTynNwx8/MO3dhm1/4RiRz8Lwlegm6OVtEEE4HejC
NJVDjqN/TgmvlrHekJz+I9e47SsjTnTfVkpOFXPlDUycCpeN5VsSxKo+DTdrtwuD
/6sPg6oheD/nAvDLQnQy2B8YlfmUvpAJnBb7S2v11XeWKi6GiuZca7TVnfe6evUn
i3JLCm/lkRc9Pt90uAPYhdpCbjrGZz69u6uwH5EMfQ04Mi2ftyyAtucpGcLufr4I
pktl5EFMEOfZ8Uc6uBFfYJhQM+tA+BlGssYFS70WUC5WQsnq1eF6wpB8kazn9byt
cEJwjXN4Y2rTN9ipSH6LF3A4VyiH0cVBymusiFtX8In6P36FRzRmuOPknbBJC0qw
5U9K7KlpU7Fq8TUdwHc4QYdWQ3cdxT3fix6TLSWJYLl85lMK7cdSocawW0sHz6hL
qzsB3OIn+qIOAmblUqkyX9kDXVQua+10YodLvLx+kNqNq3slx4z9nwEgGE5lhhpM
60fzBYOaWuwK84UnjGWDOQuKygNB8XumcJZOGnXiwO5dbdrn9yjkPN/eozcAnyak
DUTRqROOtsOc2eALFoAwKCZRfIh46f7L76PMdSQ/fx3ruFBjTGRhiciGjCM8ArHW
7MJ36aLURPOauTYFVb1m6F3h7BmsDvFRpde8LOBnh3BUM28iI3+UBlrjLDwEMF24
gGOb/IQli5cWVcImF9u+6m9KpZX/k+uCjurIL4qe/L6ZYasTeHHC4uJbAXX+BMCD
cCsZeKWyItFgfwsgtz4vIzBAb5WSfVYAWON82wPKbYWbf9dcIyvmA7gieCVQ41Gp
kRMpFQQ83HgT7zAB05+aJKXfRq6d5Ju2bU7x9wuV3lxEcWO6Lohf50nNFEZb2THr
JxTtMiihLDJk2SEqZxFcG+dy3WyIwk+1yoaEdGgm7qkEXSL2/burjpwp2UVZchui
nlV1lUUGNbPJtSE52Zp1nGUGur9lolpHSIuECF3MGH34elH60HE1g06Hb2OWq8Hu
tal+NLZoQc9nNHGpiaahPKUhLciPH22cjzyMu+KWFF5qtPWQLwu+0iJ+RM5npITv
cllIBsWbn5QVKKJUAxzQLAIo1ZuO268oZTzIJ6oDQ7pv3izDQKMbFcuoZKcElB7S
0ahw7w+IiIf6xfjknGAdKQOftEZ6Qu6yNugwFGDiL0Eg292Ba0JdiLJhkOW/WbSr
2omrODiw+n0IIj/JlHH6qyuDOxR2qZ7pUzh5g6YoOvFaPngtLCTL4Xd29o3HzhoJ
oc7S3zoMOSHxlc0Yr1kUpMCu6nT/IJ39VWM5hxvkbPI6xqQMjQP6hAWtVygA2OBQ
419IPNVmadoB6QZdz9aMwObO0EbNumSrSaO+HdBrNCFSryTIc4Ml1TU9m5W8U8rW
hD4YAinMRhG0uX8LRsZp90O9yrhp6lxf0abOYVpYPCVXrTNAtlgu6z4my1b7LXOS
omt/Z5LYI7F0l8xRXttCELgn96j9zdSBi7Bp70v4zXFsFpTNdHxiiL2ZkRoFDhAC
Mh2sRaLwOPvpAB54nw33c/uDqbUcHfwtNAw4BsCuVtl8DtEYDpPRfq+4KU0o56bF
mqzaLrXs5gCt0e4uQComn1aHRWZ7cP5KnFKpyGDrqmG/Y+MZK6bM2vqcLvCQjNys
na5VtqZxGDFc0xg2PkXssguO38HCsGKg2ODrEpZDxbq3pyTIUz61raHuAenWwupJ
GjbsRGDioVzxVz3ZUQJL5Df1cDAaayc7I++BgszHCjaMt8QtlMBGt4sXgPJyW8+G
2gSxOs3spV6kKHrNahxXyQTUrrGXco0p3RPDk2eHNYAVnR0BBxKJSAhC68DWsv4N
duSfhcSFhhIkUci8jgid7GM/vZf8YeQfQJDLK2LfG89oYQjdn0WHmphFggWiq0IC
zv+c9y0aVi6n9bPBGyzdOY0lxtus1Ul9gRwiQLwPdsjmfQxsYk9sMjOfLuWpPn68
WkNRcZRGI1JVDplKmx+KuVf1gR4hPdQiy7mpWrFlOJIu67NGKl9LIybJgq2MjIEC
jIlVsz/QI1IeXcfyc/xr632K4NS3mY7fdyxiXLMSxUfRRjEz0o2ouLXBNxr68kPz
MmfZ/LX7WBPZwIR9EN3KgVkNphbPVV81IMVHoCXcXeyJF00duQX2sNbgWUDVPk6m
/DA3rvlKwVkSlzxhxF5p4gtCCxQe/JFjRsEudBrpFBsW9HWpQSqwtMFJQjPdfyOR
hCEcZxRbB9DDlon6jW4+trgF3ECGqtYjjU6m/+o0h+T/mYaVaPuc1CPrgLyGNXpv
/l3qLYBZczyosYRh7kBj8xRqW8S8iis9th8iCnIBG/Q=
//pragma protect end_data_block
//pragma protect digest_block
tZ1VdWwKY08joXt4pNnX/0Yxjlc=
//pragma protect end_digest_block
//pragma protect end_protected
