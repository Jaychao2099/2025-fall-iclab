/**************************************************************************/
// Copyright (c) 2025, OASIS Lab
// MODULE: CONVEX
// FILE NAME: CONVEX_encrypted.v
// VERSRION: 1.0
// DATE: August 15, 2025
// AUTHOR: Chao-En Kuo, NYCU IAIS
// DESCRIPTION: ICLAB2025FALL / LAB3 / CONVEX_demo
// MODIFICATION HISTORY:
// Date                 Description
// 
/**************************************************************************/
module CONVEX
`protected
T_f5fGP<OHBPV[1Z(JI)L[=eb-4QXJCb@>;e1S1:491g4eeX]9IQ))ZO^)</c)/D
b@YB9^HC53UMZU\<T@RBZVeBD;GQ^DU)?>YC1-.DZS]\.L]Kg)^5^3KH/SR^6?)V
94QOP,@25gL6@I+_66_^SQW^6(43d4,17JQOde+/ET_BZOU-Z/NW0(Pe7;)_c87E
N]-GG4OT]?[;=S9RgePZ^2O]M8Q7C7+gN,g;[g4.A8L52[<GX+KNMGTcM=<=_NgZ
T)]BfR5K=RL5c<)\&2G+W^,8MJTfS1F0V;0LRafBVGURK\0_#O/(FIDBY7<aO-#b
fECS+5Y93@2SR_JAQ88>b#7?I/?>>d+b:[Z?B>DG.32B:YOP.AW-2M.X9<THE0Og
#MML@Og<6@-N5J\/&IUQ#=AQ1/L=IPP8GK\=N-dgBK]WR?fBcBEOS3\_1_>[cdH4
(Q-4WD.[\67B18ZM542=cd4EVD4<EMdCT;K]NgcT9R,5C=\/3K+WXde#GH:,?W=0
dQ-.,R8L1gb1/CJ,/=HU>a(1RLIEe1Yd8-;(L_>P6<5gJQ@,K3+=F@WLSafO4)W-
C#@&Eg(f[f=9#4gEG@eKV0E=[S79R:d<A)g0(9KZ@YN^L(95-ZF==B(d#7D)L?<^
QP4B\4b0[]EAFV+#<O]A1(<d18VH#?>9>E\IZ)\,cd4N_&VHVRY^[9>7YGd]@PJ_
C2WaA]e\HVTY>N3?^?+>E_5:#_NdCSQ+RBcTVfbTY4JQZ[Ba1N4gReSVOPQ=P0RK
GF+N?+e3GG4RR>D>dFHGJ,+D^</\FQ?DYc6X;XI\DgcZ&5DF,HE)YGOM?;LWD1^f
K:aJ<b::a[9D=4<JG\B]6)1A,@f)JdgCE<bb=6I.5Q-B3MPRK)7,aB.g\D\M#&10
HGZ_5M4<A_.I9?ZaHRFJ>:5:&BYJWeUf\3(\4),@^RfN1)Q7>2Zd?A9<B\d=_86)
B+fE>8^2dDF6+:Y45;CgF1;FQ<B1M&_C-_Md1J[TYGAWa=09/,e=U8T(=))VS].)
C.C?\aZ4_:GF+FX7U#S=J>;L@e_>;_&4E;gS<_8493]2H4K+BOE)Z\gD#1bH[<>Y
:<#906SHTRU@5K7Ng&T4_5J/#W:G5N+VB_\LH->@4Z0^XK_8-^2f44+1eW[5[ZW0
AMcT=M_#E>eRbUKg1(PeR&^2,E\G68;)+/17I9;3Z?P7Odb1)3)G>+X)7TIT(EBW
g#&EeNY])4=SF)4W:0WSB:-D6FVAfb42E()O+_gWTLb5@6\?87[XMYe:@U7GF3eE
Jf&F-)J\Nc528B[5CE>,KXLc[GJ4fYUA=\39\KgY\M(/#fd6fKFT4,)9<RDE0X<^
[[ECX,&FaV;KW+Wb&UD63)173G]U6bX#L>[PIPAa-RPFL3b]e]58<c0/L+c2[UcF
EGeYE-0JEUb5D;D&fS8R<2fPa;V#>IgHD,2f[;9U&>AIb_Y,WcS4Mf_d>R:B@:\7
=VU3HG.P:#IW+eAP@5&Ca)50)OaW?@)6<VL\;8OTU/H+P17PJ:#OF/TZ4KY16VN?
/Xc_K4474U?eQ#a5:fB#(&Y1d+D1X,^&6>HZGHe=NML<da3=MN4\@^SW4ZQ][Y,]
?NEJ.D0?5KV7=?B9D[QLUBPW\]BT3Z2Q4@d&4bL@1c=QJ6#dP7L8]\Gf46VB76-[
.V&@f:>/89=RQ0:-LL,<ceG7]3S7>DL@F[/\d8Mg]#0_g>FVC,TDZ,6@<C0PX;35
+U(d:4&>#L36-KVGN>TY.c87Z>_0,]OMMA0D/L133L,[L1BJHCB=If1aV)M_P\16
D>A^WLQW>^cM]W[>KOK1Ya&dQ0KNE.P=P_U]J<:E9Z9F]_QL8V9:.GKJ#Y=CI0?B
R)<#&IKF]7bYg5Yf<=)Y=BKX[>S.S;V<YGK2R8/Qg@FF:I&@/a/H_X.Q=#&F;S1S
I\E<20GU-[&^g2)4,JKH1X.Y5&Wca@dL.@I(g;7aP//_.H-(=U]b&f#g)K?fWE:-
-4)T+B@R/)fWPI#E()?7&933,e?55^C]>+A@TPNE_KfV-,Q]DJQD8J/[C?&FD+@5
LTfY>4CO_bOB75RU:>KcCKI><5.-^M=XM]aPX]_>J+_F#\#][U)_SG^EM<YVJgT7
Cf[P^85-?aDHY&RFHgQ??MFYf0T+87KH)4U6,25[OVY8?BUVRNXA7-8f<7FQ:.eE
GgN\B[&edJQ9a@-M]>/ZKZ;3MM<1AD_gV&2GLe<F-.:9^+\^V>1K2DF+&T,HGMT0
&g)EHM;)[5Be+-_@.,P132_)[5YGCg)EZS.SP1DJJ7+J.cFbF@=cZV.#L,^,,X<_
geP-^GJ\J3:QU7EYFe\NYE02+J=6B(7C_ET9FOQHRIN7DF(A9?\FQ,HVS3Z&]gW_
dMHKO]&?3:)^)+IJ/8U2\BYd?/,MJMR,gg]\A_=UQ48F?6AHJVP\A_BbLEdS2bSR
M6F-EZ?fA(EUZJ_=b#b@H)WAN_Nb1#L+D=AOLAU-cAFf3&Q=a@OH8L7HB[PE;\OS
39CX^fb]bZ[b-_c6]Y#<8ePgY)WK5d8RYS&GcKZaD?dd;943,9-XY-B/J+Z9B\23
?MWg3E:3>CIV+^1JHG2E0?B+A0^P3BK]_UPM3BKVK]]gDG3/V1gcZ&gIIN[PC=?M
dO1Z.=G^CcZG?g81QRQB.)#3+KQ3WA^e+K,CQdd>eQdg;(L;97IdR19(],Od0=)2
])6+OHP@QEYA=7-M7/g,b0BgM38\7-5+QKPN\>Ue:NQ8FS_T&W\Y1@cLD-.XgA.=
WT[],6_0L5N[90;FaW0db)DHX]>S<B=5H;?]e(@6ZXG7CACF(Z(<KV:RE&61eSB)
AZX-[,N(geTB\@(_6Q?[<[TPUNXA:HTM1MC_AL.OF><33Z].A&.:3>E:c,CdM9g:
2f1B<eB0\[2R3UbF>FRWe&OU+95T-DW.MY(#]9@;&A,9F.WKVVFY/#N1()4L=2V+
E8>g]LV[H4MgYZG6&Y1H?954YD.X7W7aJ..6X>A(d-63;WX;>@\@-P&Qb)I_ADR5
00?YVGEeaB?KfM?9:>[>B<b5:BD_&,69BgN[6:2)3bK(HT\DU4(<5&\L#:2=QZRd
]1.6H^A.d54])=[\g6?aCO<MEB,SdFFWBdHAfcPg<^?b_3JWUCK9GO#;.;R;^>;K
D=58QEb<gH9)-E(&.=M[Z5N0UUcD1Jc@T#K1<cU+\Z.M[U77XQ]^D[V@=1T\#JOZ
W<C80-,(TA+g1?cbb_eNafJK:_;F_P:7L4EC)6V7gRdGd1L=W/3N@K]YC,a=C+-F
f#_bZ8\4)X@7L1]KEb6+PHQ-#J6F-QY>>1BdL@2Z8=.H6ZZ?T#@2-,S#HVEeB@Ee
^>_:=6]<3UBdfXad(Z+&5U]--bI+YdMKY+dB>O7DTb;TKQN)]aNXFJ?2MKN(2-J?
/:f)cWN)N_7/TV)g]ZG3VafV@[RE)^86#bI[dLE>Hc,Ua1V@#MAUL>YZ4_(gO\Ff
cRJ>S]C;8AD?L_SM&LWKf82PW7NZR49&Y=gH9DM1(S<A)cO1=GKVa5LD#-#@VT<E
9=#TeE>4_NFE,=QJ)WE/@=(8VXK1UNG1=[DQX+&#4+<HaJE]1c>cYcM&0GP.@4.\
2_^[fSMce_(:YYb-BQ_Vd[;X&3B^d4&VNDQ9^8BSe<N4K&JYcSb=f/\gOT>g;JgQ
/=RP;NK6::a)]KGP#-DE7(+(4Ed2<2V7=bD@;2,_d1[;Z2BS.W,-G3YLHeV:SfDR
Q+Mc4V(/2d8DY5YM3Q_1+UgKW^200TU^^(2LCC7c82E+g[.:S(?VEZ@fFYcO_]G(
f(G0FB#6?Q3[5&ba.H02;@3W>VOKUAHEZAZ&GMB[WJPJ4b^/b7XaUSeU]+Wbb[(A
0^6JJZ<_9&MHS1L[g,UKU8A;bYW>W<+1/0JO1@[OT#B/D2[f[c_/68[_C7?Y:75c
M]bHfL(6252TRL016^WaNX)RL,b:gBF.20IaNJc0\@(>.cUC=>(0RS^4ZR&P;@-Y
R9W=g+_-/S)-R8fSFEHVL82#eHRJT&SN9OV::A6#>2L=X0c@S[SbVe@UUe./]&/P
,df_caTU[IJQI.:B1NL\BOb7O)V<DH^;f^F=ZDFRHO4cd^a^1QY]aGaB_C>H7cG;
Ob[J1^CNDO?@:N\>88]1\\-?P>][>f.ZZ5_BD\R.13Q11U?+;S<]I7T(HKgED1gF
M@3<-)P+e9(A=N&;QM?[d[83(7Z6TGUc#WDU1.N&B2Z/MF7^50<,V7bH/NX)W1ZH
_[8b36a]1H.3:(eOb7J05@:>E.I><(WeIG,2XU>-MD];=eAdQP0eUHVIK1fZZcR6
Zf#3N+S6HOVdI,H_EX1Y8R8WG&LVf429I)+&afIE.AWBf?,M2;dT:T=.Y)dO.,cI
U#g-,3<7V\/3JN>,]P_-^d,d]H_7PJ1H5g2:^0.R_@-7,CQ)R,U+BJKNeET^dd<G
Gd;_V(X.bNYJM_F=W#gQG(W\C.T@SPge_4aF;XBTBQ34=KbW:V1TO)4^ZB^,-<dS
g02X#]>6[B9<GbQYd18B8d?U5[D&\O_@(W=W-ZC^=S9XP9]H1(HR9N@9/]4=gc=8
/AXTLf7UF.QX7;J[TAQ^4_556]dBYE7+(+<g(]E&[#Q=Y5TCD]6;cfVY<FDg,7?N
[GMe.S[&/G&N@.RL_?[#/^T9:@629.M?9A5NT:KT?g_2C)#G5.WCE(f55,9(1#TA
@TO?]?HdJ:aNO+)[IRFUJ3OFQ<6SR;eA)E:\G6:3&EL+4Va=:+BD0fB&YWUX)@E4
^E3VCLVT(J)O>+_IK_WVVW2TSU4<[90/A,ZMHfO(A/>2=d\/g1CQ@@R[?9Z1I>d+
\b&6VGRPBBfFgA?ZK#S@gMEA-e9754YcNVC29T>9.e17=/(6CPDeC:ITY1[QXFX[
;^Y4BL.,,XAT-(5ZQ+TLB:T[HI62/T@,ZPF(f>2+_=cK(T6^95<QHTDTBUHAWS:0
9A4LAU9(204AD+].dQQVWU#\46/B#)9McWMAXY)3ZI_0/7JQ)?8#(H/MP(&0a#([
;2QDb9Cgf>,GK(B56b+=I(PLIFF#K9L82gLB^aLd5QFU);^2+c[c4CO21R1dGY&\
35GGO\Ua5W\B4/Zf\a(H,D?P+;2EZ:X^8)YY-A)[2W-O)5,gW/Fgb6aL?MQXOGN+
&^S^2BF9B=aa_B/@EBCWY^DC&S7@bR9PE6;a<a;M>CbVTK?\6E;F\V.=OeAcS_Ce
#g,bHQgL04=6g8\XV9VVH4<B#J6_L#WQN>7dVTL#<;,-0\-I7G/f]=[AT.^CG6N)
1RCB?9^X#V\/T)NZHF4TXL,2[D2g;DG.7Q2UY0D>&9)D.e5,gB8?0X3?38M49]@I
9fbf&+9f6;egE9,O\5D4=G/W.;D?78MQP67>C]^fcWT8S?5SP2XMJbCS#,.cCZ:6
1.06)e\+T?aXbCQ5>a^.9-NOQDJBK0M8K@<I/9_>QS^6U@M1TdCWT8@PHI2],,:-
XOa_d,S+Z&S,IF:>69:.TND-:<VEG8AT0a(I3_FP1O2AFa)44-?ZfF[UIgT?Mg]8
-JW3M-GM_?8)e>B]<HC4K\V_d3=<-Y:d93]35G(1XGX(d;T^a;[2>P]gf:>DG^X7
>7P9Dce_aSbcF1N7B4+-0#?<cJ];IPH/K^PXJ60&PMbIC5N=TQMb?Ob1_9SVRdY-
gLCHS02O0C=LbUgBETdW=@Y9Pb(4G>e-L.U(RI\^>1B6d4:eKIEQ,>R-(S/C^0\(
FAAB++J)NV+X/f^+1\69TYd(f7ba5YVCgS<DUJN(5BSJ(PPfJGc@AgUXfOZQ34]R
3O5YDM-NQ3f)Va)Z\NRUU(/J5f#8XU8DaJ./BeEIHI@eQA-I6aYG/YUfHLK?F2b4
aKR1#9O7_B\HAK@eK47eLD<TP6R]9a8MQCAbGV[f?2:Y:&eM^6)9I1-D52EQ7K1&
&Ye<aJdK.ePfXRUAY+H>Ra,WOTb,-E+beeHQNb384MS^HTTa_(,O+1>U]I)P@aXD
8VHOOH1c2HVOITg&WV[c^??<?f=5\KM)0+Z4fB:F7#>YZ3ITgeUOf;3gb,@A,f9D
=b:@0cb4SN5c8:g=f3KK)Z1([.^2&:(F_]1BK9&3DCcD_CR4/b(E:I/,[8[=fBbL
<A[53)/^JfL<8_Z\9[MRWDO9eL]<Y.(TU;0CGJcaTfWI06#E57_7]BAK4#._&5gQ
^T9(/O.2&3QRU7S7aGIYG1:F#W=D2JDMR+^M5gNa=#W2Pa#He)P[]^IBIX]LL&3=
cBBc1/RCXZ&9JJN)BQ(=VD5><Pd[&ADXPe4ecYH81VHTTIbLV8-7#E;^XA__)f?+
2gY6ULZ)K5^=DOL85d&I2Q)FB=R&\eSVCT@S:0MYNf6EY:_WV0d.eBb>INHDgQ)]
R1+7dIG=BSE\5eEX7d_)NG-Y>@D8J,9,fEKMBI&,;XTZPF8=JA7T;7bU_Vd><DfB
d>GXW-87-FU/2VKC])bc5X=a.[dI\_[):+U7ZbR4@Q>9+4M+(6bCLgS.J03QWB_T
=,T/d#M7_J8HSQ^M/,2^F1RRF1?<eQC:aFcZYb0=\LDecSPL:=91d;T?MA>Z<FAf
7J(I(&<eg;P\dDSWZ(W\6Hff/C;#XbdagZT,.b^8&]eA>c0aLPUaP2#5;7Fa.VN,
AJ);2=cCES31RWSCM629(J,J&4Ng\3ONXQQ2/,Sa3IRc0/0AacR#[dGZWY.V/3+P
M<#=QJTS.&A8(UJ88ZE9(>SS1EPU]MMEEaUOY_AFY?>=J<4WI.OY8XQ(2O#3BAHB
2@B/>?::Qd49F,9=Td9W<4YZG=CD<FCBW;b._/A<SVXP,]+370GLeKYL&GC5ET&?
J/Y1ZU2e[HT4Ve(3HN88CGEe#Ua)bZQ3:e3LI9V-T=8cS/,9g[YG:fA[SY#1CFN\
M[/8d8VTX.=+1f5XX:aZHRa]g+6HO3]C60UG30&@H5,Y3GH;g;Q9EO[?EScRX/TW
c5RM+g8];X7)C?BE/S?EA9c/WX/^UKeDF74b?_WI01I).3,4fT_--b6&:U<[<WRF
aU=MY]W\R_B0SF]Wf9<O&SS>-GCP#:fLEFA7O\eaM)+W9Z4\JeJfE?2Kd3^dBg82
4=4?4E7E-fZQNE-MAeVE_ABTVF9>HP0?M6\>O)FeI7GZ+2]4NRUCV6>:\T;:CfL<
2E=Q9\12dW?)dOI6ZV<X?bbWDO&\)DM36S6)7R3>UcPMH/=5aKK]A#-b]R2/Sf8[
#M<g(8<(05X(B<5<Db_E?\(3##C[d78]=5^8?:1QZLBbQLOQ27aGV[2J\N[O4-A;
2:\#)8NBGEJHDM.8EN]_D>A>NeeDI&EZCG]I^JYW-^cN1Q>4FWVJ?LC?+YSLOef\
VbLO4M/&;aCWQ@F4X(^1O.R9YZc/dTT^\=6JT3>QOfgG.2BRR90UY&Peg(DQF.FP
JPg\\&NP<=a&P8bYV>C2KCcZ^RA&I=g7ae&XU5=f,-I9I-C4_,<T3G]68D^D2G.-
c4?,2#a<c6e7M8JbZbaZJ)+6FNKK_;CdL;7KLQ.Da09aXVXRDCOOWb\b\Z]XR5>V
@(feO0(1J^U(d4c9-Oe5U66#CSYGUA[fBRDcMFQ-\QgD2\ST[<4RLNI\]Ng(FJY(
]T@+.\e+2)42YJ/#J\aW]g\Wgag/NH/G\2\?CWDM6?4S0a]/JAPc@4L+81,.S9bE
):ac?><@I0(Z_C8--B,CJ.URI_X8aU>2[g3)LaKJR]AA#b&<A_3N;M1<Bc5eF:JA
X<CXDSL<52Z@><<6LD/4F-.MfO=I4KS-0T?=;VM3P0_9Tg4]8YPWUH_4)e/E1:N]
#gPRYgJC0gAE8^b0?JUU0V]TP](bKg90GMK5906a(;QNF;W?IPQMK(X\X@LULf:3
SF<gS7?BTG(FSYN/INLa5?M&(66d_N=:?L]A:DacSc2OC(+AHbK<VGO#Lc+VU>LE
PS#O1REQ+;>P.AXY2cCXS6(;@>)A9G;d6eT#17g5ZN\W;.P-_PMf.-IJ><a<)F8R
Cd\M.K[0(A9B];0I.?c)G;)0a+S^J&VbP)6:]QCNY]SDGG8,eDQXX+5BGf\+G#_)
]Eg<QYXP6WfWgaDRLGfS,\(Q^<<]B^>W>NJA9<)=/a86=R+:(db&3Xc;Z:#A\T(-
<>3<:GfLa()a5;D(bVFUBAL(c3E(?2.M&])fL@^]VU3+@[Ic&f-)VHB/#77-&X7(
d;YQS9RaA#&:da-0KKcWd]eY4I9O_OY1;Ve,B4aX8CY+L.[.PRX=]-0#AX??SDZY
a?,?>GW@SZ5[1<G5.@g0e@Aa6:H:CS7P-#6I,YO-Hgg>&;95R\T/dIDOOZc]+<:>
)K/&7#2[:@?agU(/+.4BO#c?(QEKJ)b),J>8M,#2eS]Ke?-3,I+KcF?@PYK0Ag@@
3]Fd>=d0@RGDDgB1N\ULU6Y@]];_.geSLIJ5CE0YUF>9bg\Xa_R25c6GNgF]N;.(
0<87:]-&,Oe^)LP?-]T+SB#F+S;2V=U\7\((_aUSXN,>2J,=RC[^c=bb-JITZY7L
UY_Z,P?GYa@#-527])G<P51<JPK?Y=\He.<C_K7c9R7gBEV@\<efZ8T_ff=T;cX_
SbO(1_,(QTNTOOX>Yf4DI8IZRAbZD57U8J4Gg8V&V/TFgVKDWDO#X<fLWT10S-dZ
[\;T4d3[eV=OB8?5D/W5NdC@<P>Y7\UWg7SXL9ZZ7AXI5=C3,-&<M>DIKW():VLX
J0Nd?3M]HQ(6D15MB=E]0RZH0^#EGeMD82PcS]f44K(^?X9MafO5KX75N;We0/7:
W),4L[\N?ET=64+W.cD&_IK.^]f-EbPJKTH33S=3H^6GeP,<TN^/QO8O@3JAe>Gg
;TSL@ZG5fe2@M/55V?O=?]G0BMN_-MYWBA>=JV@e5AIAV=^[aF._9^F40.3_JXS)
IB)OYf&L?\-\=?LQXfcWce]70f0172<P6LEeQ8BHFR1BWbaO;f@6/ZSE4.VQEJ_;
,H+g;.W]-a?&,J+KeZPP\MM94)@7>e:K9G[E_?Y\TW<@.RPa.N#C2U51MfD9-OT8
b_cT+NTDScX4T&eHKU,561\PK:+A#ZW8]:7c#U@X,L=V+GMB82;f&RQ3E;PIW#g=
5bLLNS8(CQ<TK<;\IE,cDd@EgY9&OfdL\:Y7E+Q^_DZZE[4:3f^b&R;OHG4.5H53
\FP3\b4_R-FggN=IXU/ON8bD8>FZI+f1ZaPQ7ZT05E6V\+6-@AU(N&g92G4\TE6I
:VSJfLKOab0_Q4:6>]:Of4Oc(f.Z(GZNSV4&dDT17I3Kg5NG^-PQ)TU-P9a<b\#H
E9L/_MA))7HPWc=3OZRE?US@+ZWVf(T=E]H4-<GU^46.WQ++[4[)2bIG\P>DeFed
\FeVLeLWD3_0.:Ma1?Q1VZ27SIBG_Bc#S+GC4..NcM;G[:Fae9aG[CH6^&MSM=?;
bGXX)aIXH9QTfHUW;[LW#X8M7J>LZ)#BVfW82JA2&GF1_\P&)59d[TgJ40b8.N1e
EeS1)Da-RJAKbJ&OTb1dW_)NO.81\7U\N=/QHIN(X.Bb=\Fd#6_)5[7Ta<09M7O/
BF^T\STZK5E#B)NJEf4KQ.gJ[-+[\=\b]U_V3G39:C4(PHK9A)XM.WLcTePMLe2=
<KH29b-G4BRb_;RF#2,ZfAVKVPVYbb_7G+C(P]B#gQO.ATAIRST2QE-#V-\SX:[T
cFU,Cd:E8Q-TG,3=gX587-S]bY8Z>&?Z<?P5OaL)-G.SQGL=#58..^T<7W)=7@NA
GY&#2[K3,.H;O&\;[>6[J(2D#[XgJK_D#T._+=3I^R&AJ5?@/,+>@f#)]FBL^E)K
_>41(WE#U(P8HXS#V?g.O@,]DX3&X.4XDS5>FI@;;b=g1.MF;=c>UEITdGXSFbPT
U8<&=aR2F;#U(U;R&J^9:a\aZC1BV9BfU?GfbEE)aC1:Kf/G/>CIC\(C^YB&@.2Q
++81HN7M:E3Z;3ZWDbaV#3S(M1B2LEd?TLc7gd1QXQSW&7SE?LZW<H?0:S<([BJb
:EZ,&1Y-[5-J?^Q41cIJV?F(S>O6B-,Jg#CZ&6eZRac.@(#[6\-##@f:B:f7>O0F
g77MP>f=&bH/geJ_YBQ[6Sa#9eXg<gU\Z+>BcD:K7@;G2gB5ER1cTPbAZD8,4M-&
S^W/],75EI9<Q6b=+?IU1BP6c:<WN)/\OU/e.G]J<S,\H[0)ZL09gXKVU,=;4>e#
&8Z19^_S#9_X1:,F=b#;&Xc8KB>,W1FMRd<6K<C?:A61>3QLASDIOX-_[PUZ(<Z7
.Ef#IC)<<ZG[F\WPXaCe@1@_caB-LO-0\fS&#R:M>/M=[I<,=g8SD.?dc@I,>VRY
1X7Q+XD2Y@WJELDWX<>7<>;6NMEA12Nd7V?<FbHIH5T:I4=2)?A8=]OHV+_CC9_5
E6W[VC&.R/)6f^M/68@SJKIP7/(L6dP3K_Z1TXfHS9LNBe4HHJM=B>a3-I.:MTP0
QLc,,8f/+]^9/G:^57)+2_0O0,YY3KL47&BJJN0.709@PW.#;-=_f]I?S:Z4BW52
\eSOc]_V#7YV<N;Seg[dY11JR(LgO<7SfRKGV>R58>@1R80]U)L^^FgZa&+JgW2S
QC+8K.J5YX/cc+U6C@F#2M.:;#<,Hf6&0HNTg5\Q#Z:Od1:&X8@f+4SaO#b5EEgR
9N1DD8PV^cUMTe69YP&OIG-:CR8S(7&IRAT4S6++eCJ-F2>&<6R,WgR+g1OWL(F2
C]+/H2]5cT7O0,gI,A5.Y>4NJ>5V&LT4cI)fAJf3KJ1)f:WEZFCJWI4H(&9>0LSO
]BR:^;C7D3]:&a575>_#Jaf\D^@c1V_5QeM(N1GaF88]#.@.C9de_F(2Od_28,E[
7&Y4RIIE8L18-3ZXLSC>aE^Cac-L/YW2<da:],>VQ9U8>W/c_444H81&eEY6C8+R
#Vb;[,UT\d#Q;..5AX\7[@.W_Cbe9]M^V)1&[\b\2I#Rf3I-N4.Q>?FJ<OS11DM\
f&<Jf7:X2Q]_8[&+eYY=F]\MGVTL7WR;c#,;&=</.1O<,;f[U_F.(f_8(@]4H&,#
66X4:.?FP1V[).6-<Hf:T-cNY]5Uf>If=Y8WYS0];KCKM]Z8(;Y>[46JHI-+T);K
aV,1@B07)SedR\EYFfG9@^Ab]Pe(@QCB@B;307Sf[[R67U32begLJ5UYcQJJ?X/,
1QH>+C,\R.Xf>B3_O&b@A<P((#:[7L(9\I]=;BF;)XXV]3P_(;,34L(e;T0.JZ=R
)EM4^;Q[I=_/dGM>cI(8D4(:8=]7[..6T/D79a?4L-L2^<>SDa5e=GRR+0=Jd;dQ
&,5ebHU#FLFJV2:2>g4S+,)16W5_f-#2V(-+eU41)2W[Z2I-aC=N,9_\?E]:315Y
g.X8H2_G91N65D3fX\7KD)8MAeKP?KU=dB5&EJdK\f5E-2_A.Y(>/)La76K<PPS1
d3A2QCVTWAT11?XZBReJ[&P5X\-1&Q0@ALJ>[bJB<aJQLL_\.HUgLO3bBRe.ZW4/
<8>KEAgGEX.9=Da/45;ANP8(edWO-W=>4O@(^(/7Ig0DJP5K&H4_7[G[AcCXO2bO
BUUY58^IMa\8(aXcJ->,XLe+0OU5[(7-)2SG0E>T&cb=8&&/Y^0BHHQ8OfH(;:3.
S;^C_V-I]&1[0_/CT_QGY&[B/[1S4N=BZcN9(OKWBRdXL0X[\Z#_g7FK7&7.J[=>
U\?8HgX_10=PR^U79:T=Y<8OfW9E7\(N\L0g\Z?U.D@[d81GKLW6G+YZ6[d\EBL3
O]K91d339]+L.8g7G[bSF#-cXS3):/(O-AW2T\]e8@?]SI>G>4(XQdVL;TbKeG8F
8Y1F.Z;H6&;??D3Ke=cg,<0H0#E(;GHE6,.),^c)Jg9NfX<L<H8^R>L,4e;V^R2+
g</Y1R^4<S5@XL6T]0KG3b5\I?d^VVd-d#Wb?M\7,D;U\Rbf8TBLD+(Y@SX4<<VD
/;>0#?f;W4g^6SO:(ZWGKQ/0cfQa3M#_f:]f5(a;\<H>NKAgXFJB,TF?\^;2Y[Kd
F7I)9ZYY-9dO,^4e8-@cO+Z^8&cM2\GF+[J6QWXa?g+?7^bOTOUP4K^+./[I[<>-
6U97.W,b,^LMNB-WR.ZaXM8d\PD/3Y=-5=NUGFLG3JTYTXa=:1-2TMea9(F)2J-+
PRcBaY#P[S2?fb_B=J#<9I_]HD]83<[F[HJ_-ON]WR5SXfH\^R2&_Q]535R+XAcP
QU/2,K\(9S;9^8RKM+YX-17T#K\U2Cf<VP=5:f#N+X[:@7ZAOQ=(W):K(PMGW9.>
L1291OK29]>DUVZQOF^c?0&OJb6aLKH/#WJ/N&Y]V5:Y8b]=f4L_F[&JM:21)daI
N0C,WVV-[7&:g#F1]6TCJDC5W(5_9[0ZD<>,^&D7&2TeGdJ0K]U6)RV>1@[N(,5#
#f+2g:U=&BUUA&_S3+4Bff-5]_=(eV_L<S\C6g:K+Qe3\Jb:?=YJ(NC&Bdeb7K(J
^>6bY6@NIPKW;DMZ9+J1>_R&-H&>=O-F=EBWCFV6L6RbGH6,0#?aWV.LRf=_TBUC
XTY)N#4;R+gbe_(;E#B^L=BDcSg#I989ZeB+b/.COO+_3;.YOD6X+)C@25WV#g67
SGRGM<ZX#+W)X[W=g#O>L]&@HWJEKGaYG#T3Q7#=&)RKad05G0BA4gMaKY\#3,0<
8a#d806e>P_58F0b(MIJ6[M<HV5FAPRQAYP4A5T477fDUA+cd&&W5<Td:1:BdWDK
#@)>;ZQKLgA+a1aT^[aP&+CK\H//5^K3Db+4E+;NOMZW55b_8+5D[B(6eU<Rd+L?
6V^]ARGM\#&&4TA_[\RG6gE#I)dO/M@];L3IL]H9L^bN.GYDRGEfSd(6f/R8-A]c
(IYERI=QFMB<#&AS?WbT#OVS,:.TV>I:\9C[E/O>4KXR78^Q_U<B)<L:2K6VC)KB
?EZ3-agO\<.)GF#g2&AdY7BddfadWPeSJ:M\>/K\LNO16Rc9QO>?0EcWA;]L=d;8
25#]>4K@JX_/S\C]4@LUPQJOF4cJ)UUBYG\R<U6(U<B@PWX9[-AKWF#\aY//]7&e
4<\0_38+S)>,-DR[>AL,^LEYa6<A)HN^+=N15Y-^1SG(?>9A/#\B&O0a=M4K>2LC
AE./DfBBBT]5<H1eLT7#VbcHRQ>a6D<?Bg15\-23<A]95#Jg#<Xd31PV;fB\#\VP
?VW\Ebe7\3(Ie:[-^?+c3O+3@fW1]g@3):SO2PK8RUYg:G2U)0[JIbYS;gOc;O9B
FddA@Gd7+;V1+D-W]fE.75=&)Y/PXe@\[WS>,#6[J.I8bBI;BZ]=,f3>7(U#G9O(
D]<&-(7S:)d9-./)H)FcDR5TP7DM)OaA4ASLbJf0^VRb:eEE[6Ua0(5If(e3R@A^
)2#?6J<5AM:17bb&e^37VA3VF[Q-T>R:M3KSFTIWI--ABd)03c\&.W8K,9(HLBS]
.MdPaR-2fKN&@RVg@2IS\fP#X4BWMH28<a2#>5R55,>U12]a9gIcI88:<WZ?2eU\
]5+.23G@8aPC[)+(>74+V#R7JK1LD0#F,afYD5Y#W<=:WI>O.MEb.McbffGQX\>=
D7f,OFBFGe>I=G=67A3-_)8=a<[M)06C\F;De]e.FJ5ZOZQDNEbaZUPGU:8MCO_g
[HC3[WS=>V?Og,1176Y;U#]WKCc2d0eL@]&Z[-+SfNL+.)K?W164EUfQMJ9S??)N
&_ZX\)cO9AVeabfTB;4=JJEJ8YDZ@0[A4d;<[Gef=eKQ.6(C-N6[B85e#_;R^c5&
6ZKMZ&bc\@TQJGe^QMY,)FEAW1@0bUE1=-VHVe)@[,>)LdY5a4bc7GedWY:P_I@U
Q69J_EJ#S[8_8[:aK.^A77b,F(IQ[6QaXc4/]35.(&7MLYb)+<G&84gg9W@_]3Zb
GNFJ(S+bAYc)<8,;W\>=UZS+FNQP)@eSHfB=SfA5P2&5c(1_UOV,bZXBcb8DYOb4
;8LKV?JDL.b,;=4X<O;4S@<[,AdY96#Y+SH0H+JB&\\1UW8&>LNF[a&\PIX4,B^7
XE(J#DEH)@M8gYA);.#23I.=K0_S4:c#=>7^gZbH1](SF0QB#,LH0^1Mcb]J](PS
+Oe9(AVS.A:LGe@+g<D#90HLAK]a@,-M-fZVXAV>5)(1^^/;PM>BFQ5BYR7W+LO]
G9O.;NE,<6IM76<_839g[f<<,+3UE=0D9^0BD.065Pdc;Q&AHeaY&35(-UO/f&NP
3.\[ceO<]-7I(>bEC8R9B?\D_W\8cZ<ce0GfYR=A;@I;\.6^;O/-U,NMb?8.U)I5
J/FCMS05LL[9ULeONK\K+c+LI5[UN4:5)P>E[+(Ae-aZ>FN(+)0:S9(L>9&RAD]0
0^MR&>ZKR0\SbP<[gA(?9U7Q=VQOYY#O\ZDZ_#:Y#^c(QW(0Z2b;?9I&C(cY]X+V
&+#SOAaHP?Kf]e?U:.,CN=5(^aS[?L3Q+#[WM;g#;4&3NB>=fPR+ZVc0_Q@JSKEE
H<FW;69fHX>-CA>^FKA))J4,6X<C?ZX&E7T,UR4N.3Cfde;aP+2c<Tb?aWeXDTT+
95ZcSdMMO8&=dGEA,,K124bc+OVTEVc?dD=_.a/VBCafS\6(>bW[YRL.6PPJ>W,,
442=^2U2#>af8=D8QLKfEeT^+]Y)V2H6<D<U39B2@R.8+?(I[((6=5c.#A&W<JFS
>:YC3fOB-T]E:TOd_ND<R<2VLL0cOcSH<37dBRD8Y+5O&>;(#G&0XdTH;O-@=WW2
W0gZL\(eI2^]R@MY/-=3g?4Ee99_fWJ:G.>9Z\J5)F34f8)]_R,3bZRAHcCVf5RQ
^Id:S>.0PD#9OVcICS=4;B49>I^_:Z[[a:@WJ]Y/566eW.68OLI/,#K9^c-UeIV-
Y,645<ZeO=S]DU^,CMUFQDW\[Y3&^T(b1(JLEETL2=&VTT.\c1<<a?Y.b:_T81O<
:1Zff?[;9GBYB@3f&KO/M3cKcg8I?^-(\WC<Q.^H,eF,-OH[B-W+DQ0@#)7D(WO/
Zg4I(IR4/93&N61Z#>Pd2)=aa6UbCFDD._P88,0AKFMM1a@?6H8G&Za5G[A[K/?@
I#S:dKcHed)PKf[H+GJ5_TEe)\R#=D4/SM&=:cW&c:d(,W)8S8=QBV]#.0@LB.@(
T71aEW00:O9CSF6=\G9_R][J(f^]IN+ZCRGFNJD&KH=6EA,873>Ie?5N>W&=6,&H
JdR&5Q)fb+S10;CTbQET+F1;>4G>AB9#U#+HAaZb0KE<YB48B@Rg[)F[))g?F4Z4
O2CAJ?(CA[=(eb#Z#@C8Z(^Jc&76B#)C\GfBM<HFXg9T7(.a@1?8F;XOT)?98:03
\\K[TWTN+9gO.I_c,RZ2<2.H>OcU+K4ZD>EcOA24Q]7(^>GP5>8E1bU:aTfBI64E
_)CaHG:S6[7.Q&IBK,MJ>+3AOQY1TEL2gRKOEC]DQ;-c)-AR@\ICJJ8PI3K=.H>a
d3>]1:&?AV-WY=5R7C/LY47>-CceSU^8A#VegBTXZ3CN@2&eLBGU4:A6M4^3M8(X
@?48R[)f>M-9eEUY-.e0D=O;3_#^WX65+=F>8[]\bI28SGJ9RKIPSJ0@?4<U#]-&
aPB<^6=(E36LCLF<X4fIK^MY\+cKda1WB5FKX?]Z]Y2&2fLS81TM]HA6aQ]5KV03
Q@A,[5^3&bTfGR[YZ-IDQ4+/J;++(:D]&;-Fg?DEZ:ZM93eG3RF-/#N2cU\J49=C
\Bac]>(^8UJX]H\X+MC#3^XJAP]YIPO,(^L\43=D6;Yc[/g2\ca+,/4XcYSH>F+5
-RU;7.+QZ]\K8_=[GI1a)Ja:\4JfQ3XTRfC([JLFY@(Ib8UXJ-:DL\DX)K(ReZDX
31;YRc&#;ZZf;+P95^X.6[Z(_D:2Hbd)YJR=9]6Z+Y\4OdCQNTI/\e4A2RTR[[+S
dDTLS0IW[b)3A>;,4(UZ07X&a_-7&-4LSF4<?ZM,eNPgfgK(HE)/CTER:[3</K/?
<g&+K,)KSHN#_^HCI)K\,;]N+KDGQ.5#I(b13.,WTRf#a#X/Z/3SW()D/47,NMA.
;4Cg,+LPTPVc&dBWf2H_0fc@QWT]\U_JBN;Kg]#ZV>U.g/R95fTDKO+9[ZG061-,
WIL.<Le3LS>8VZMg)e\e/9e#AMLO@U[6]GNgcRa=g@8W>2R__fdB>)Z0fbR3.MQ,
I808^>3>PF?cU(D2IDO4L\6_W,K8eHTO7>3N88_;;7OD-0,L9X[gMBMP_+=6XJ]L
b@dS;P77Z1G&JFVQ;XR))3DXEKb#VA+7g.P8M1G@(d?.Ib>,</eDD^:AO,&?0IWW
J^@UOT2[4987UWGK9937IVWLZZJ\H+&ad/?/J4R,J/,cBQM?N31/9b#2N19BT(66
]-G&e@cO.@DL+8#H2+03KfU#6QA-c79XE31M#/YQ5H0Z5^/abNS8R[@d/+aD7218
fO2..K-@+2=]QJ(JNP+bQWTDW1Y]?,W[XE&Fc@7)V_fRF8KE@J#G-USE#]T0+79/
a#D#Qd]&KN9eGD@<D).1ZJ^DdDJV[;64XQ:-_M+E#6IFGWaHe6_#_XY?24)/W,,M
6bD,P8ZM5A:U_e4A:D3DS(R^8eKO@RS-[7aP)/U@IVQ>YMK2J2dWAGIBG#^&5EOJ
:[.1VV7K6L=6A4-3dbQ5F<ECQ>RDJ^J6^b^XR<_V30M:EF>NHYB,^edN(@UCL,W4
#a68@]@-a]4VR=ZWH1XDecK_ON#1ET\U:\gIB](GTANdZO\\?X5A=@4N)_d3eDMA
5HY=KEcD(H.GIR_5JFMaR\EU>a&M7B1N/RXA/OVfDbV>]RWe0=F?;4HbPW__Pg@c
9Ie>:/J]:Z&:5Ua;PA&g0:HB;3\W(,0<<XU:/<.,]TEX<\3BL:0)bT^U.E4SD[+V
<d?2^T0_ZQMXH\b/CV(-LT(3CSJJbZ?RSHI#b.>3[F/X8?M6+RR?-R.;:FMWD[F1
H>?@OD?LK<^g[53.XLc@e/>5D[d(UW6?3&4gV#.Qc&E_?N&:B_(XE_>FF/&@)H3;
3@=X-M+(L(5,S)6<&F:B<Zac-KNHZPAY+(VE?UTQPVYI4.5K^6>F0G9A(dLLJ=#[
[&-CDT23D[NU:1QTB^3R[bB&C-K\McgRGACRV,D^=E.:OII73gLUX9Z/O/+0OVd(
PC5H=#cFFY;L_E8Z+g0?ZG954Z,9Ze7aKLcIgg(=35W+78@TcDRSIA=5QRZ&X-Q:
S+=:>DB)e8QbF3/?&##eBDLIC@00e5E:WSJ-L=B7Q0EE57R<&;F)2GTA<\8WVNaf
Y()-MF#fI0(Fa^0(+@XXX;ZZFP[[)@4:R^^_eM7+?GOJKKQBZQf^8bMdJ-eRU&Z:
PC[@[BTO5fH018[fWI(e.:Y1=@gU1129UY<S[2FP3]6,A.:JFYC2#IeNPC>=P-Fe
U91IQCB0,J?8RY-WT/G/@A>7P>Z>aX]-(3=S_@M976YUU/L45d_4b8_3PT22Ya^I
X68f;Y==)[?5Z#>^<a_VQ&JMB2M5OLAY&0d02Z3FA8H\::TC]N)2#UfX>?gW>^bW
7eB666)J,b]U51)U+SWG_-3Pe4K\E/(5Q[N23)/=KH@D=:<6cH8/<K;K>D3@TGOJ
:_36,F;S-CUca&;agT-Y=F34dR9f8YE>\7aER\JEO^_K3[(,-gC[J2&R(cdAQR2T
B)L-;T]4<2<FAE9=]aFCD@WCgOS1Z+gZ(g[DD-fGF9QNJ>6V9&+O;CQ.TK/J985^
D+(g6-7WHdfCgXR@?^:b+5+Y5LDI-9,F\R+YTcZ]bH[9aX1?)@>./>\PH.A)6]eC
N-K@KD_L88AW3FRAEZA<OMf7B+ZS?FS\)ea9J9&aS#FWDcV,C)bJO5Nc&\A0BED1
R@H.8U=:N_1BY7gB@fE^/A#a[S[MZP3&D>^3A4[UMJU4S?R^.?[gGXFLaEY8WgRG
f>E3[KC1Og4:CcE8P[-ObL[:TEaFD@;c/C\^EYRARXK)e\&AUR+^SD3RM#CJOe]d
<4]]ARVeUPb>2Ne,9Rg6CX-d\PJ3V@I3=#\-TB/#SGH:R0>7IW0CXMQX;2)&FONW
-DS,;5f4_e_RJcN^2C>CJYMW=6YaG6e3N9+BAR06fR;W;9G/G+RUIU>GJERJAJ=/
1[7Gd[Ff;PI:DD&@A(3OZ8Q#@=Q>80A-G)@XVWb?d].?Fb]F64dB9-ZWL&CKAADG
KOW#UGXGI5Q]=DEI,HIbD[CC+2VJOUQ(H4fge9F,7D2R_a+EX)8LU#B-)M4>cVDT
[/D45d8SVI8\#b7Ra+0ODU#D5]P9\ACVJ3DRBAKK;[8Z4Hg@MMe2A)RNB\##d))a
f>_\OH5,MTW>]=V:CD+]9XZI^>SGGRX4A\N,5LPAa;Z#bOD8-L694KZDP/33ceW+
1Oc1[\=Ca8DIPGMI89/G745@eM)8.L5/[)-G\K7W1/28,^#,V98NP#1]?Q4[Fd3(
dD&?P(Mg7JG)P\B6>,&2L2>gA>OV\;&>BEC=XR^M]\2L:.bRQPJeB+.1DH5T[Rd.
1a2]<3_>=,^=bWQ-OO55H2e?B)eO\W4abHHd3=Z/W]U,4OZIK)dF&S5^Z62\Y:I5
\B?N4Nec9XGZ\USWgNS01BD?:<Y7Hg??M.T5;07<<13U[dB1T^&_?YB&&E=La=^5
@ZZDe_X@;QbY9cCJRE88W(2cHe057@aXgA+AL.E]=SeBQEG8LY?=Ag]E<U^6VK^U
>J?B26H>a8;2gI6f/G:7^Y6H+U6\bR34?<b1[R+NG<;,W9^=PW,P;5A;N..E^9N#
NDc:JHOO;)=JH6E1FaMCFIe&HT]]:cEC=ef)>#N42KR2Z[N]5-:/G=9HD#E4Ve[(
0@Ra0+JY3NV/V9IM_4GELN.d?>IC/5K_)FT9,[S?+[\/P5f4C.R3JC-1d/e1VKBE
b;P3O3\==QT^Y[d0aBIIa;BN=F7N:RF[MeJRd9g7,=G\SS/7];D=UQ/>,TI0e82[
P,97R\_E,D7ggbW41HKL3-,#V0f_[SBQ:U83VB5)BBAQ5/3-/deSQYcV[^g-C:)M
2T-\U5K?&Q]7F<TLAA[X@fPVFP6D(CU-<>[V?dfaJKO0O#))B1?HQ#,ZGP2aJ8>A
R<XJfVaMFP#f\17gKGF9E6>OV;4S-d7@+Wa54.49>N?;XLeI7__2-,g+FE_bHZ9V
TIcbE-XM#ZJ>I^fKaK/HRdGd#J,2+E;DTMHK>,;;Y6D9BO=J[P7@dFOLXSPDTGV]
+<2<EQgB13Y)6eU3gFRIK<ea#_e-G/f_6L)OD#0]G.-X;eK0aB\:)D#O4LW&]\LL
0T0:[/_2dWXINL1NEEC^X@ebGL&AZD7J?(3]BZ.52.1]#\0U.FF9E_JX6-\I:>1C
W,7NR=DF&[_F(@b@J(g##=]Z(#T4002>T(eM1d(^cF9)Z?Fe&a<Ld_84;-#7AFW?
,3J50>4_9WYLW>W3BX?YDCJN^A\bM1f77-8H0=d2EQa_R?d@X3cG[(9CW2\b7)?1
0W6KC3aP=0#.,I5IB,NQ41eXZ0cFTc@WR9M_?d&9U]cLKI/6\+ZEA125=.GKg+IR
KA#L)C^(Wd3<2b#F:>1(MJ<M@?6AM3R_UNfV66e5Tb.:gC29\/W84b)#c.R40_c)
@5N9TWJ?\Y66V,ZaB<fDdUQ\4gE=[9.(AZZ-K4<W5@X\8<9AaMZ_MF]Qe:R.YaKI
,5bJCP1<LFUM4V[&bTKgB_\aRLEHG.T_EFcH3;867Q\\O0:2(afCgXa[<Y3eeXFb
[?7FcKbcLHe?#&:<+QRO[\;IL[a(JCMQ+#:2/S0ITNCa\?Hd0+0QR)7ACb?2\1AI
?MU@-SU\Na0=4aGC@4@H.V_>gc>>VC2P1BU>R+W:?@Q<0&MDGV#_=UVT[O/?\\c/
8@d18)/+NV[+3FO3V]KV-URS4-a]gZgdaT/Zcb\#.]Qe]N31YNC)@X/FG19d3^(X
O5aS(I9VfYgb<=Rc/L2S1.GcQ0ec6/QEY0:N+5M\\eVN;_W:8\:E+cf+.M17_63[
7]9CY_B;[3_OQ3;BJLgc;B3Z^-^G@2TLD./&>.6R>LCe8PI=QP1d(J8]>A2QU-Ce
c3WELG>AINagF,f-+[F;&K[WL>)e+JRW=Me6-+BULgS/0X?YbKMD&-B9C5IMLCX&
7ZJe)U)<8\1+G@]#<4,PIFeS@dW66H,1/KSg.K#MEO=AN01Jg.efO4+Q@3c>::(F
F?@;I6A0HeGZMRdOIRXMO)E5:-<Q<THd^8(NU49X]27AG$
`endprotected
endmodule

module SUBMODULE_1
`protected
?D9gNVP#2JX=2EVFBVf6-55-WD\+Ib,\5I-0KP.6(,)&SGLXK&;^3)MaPG;_&VH,
K)O>UN9g3^S\&eHT#3^6IH:Ua9Bg@;394cJ3<[\E<1[TLA&FKTXL7&aR.U0Q82-.
]g#^NEWKNAe/_=IUOG=gEb\5,NggA>@bE8R_MKG9]#\,4>F4CJ>,G^I_M,ZXDCS7
(;4LA:DG<?<H(dZ\cdS^D(?EI?UE+cXO3>69TP+.@4FHKJg66RU<=5cTFd@_4(Ia
E>^DP/eM02/(\:d;)FLU<_-cO[_db99QMA>e-<FF<KNJfT>egd/I@DXY-:[._V:Q
H\6?N^Z1[-C.58d_dK/6K/^6ZVD[6#,P0W#>,&P]_0>7Tg,9;E(O@CbH^b>IYW4_
dQI481[5@BTZNgBEJWAU(41?e+c&FZVOLPQKd)^R)JV>R=ORF2EJP:E_ANe4[OKS
G-QM:;ZC\>a4d5a<,LW(U8D=9gdJ>5DI&]-SeDQd@KJRG(4KQbV:a^.(3^>C^c5U
D)7HG-fV?&7g.eLe95W[KJ;K)-aC>F@M0.VD^\NaTB67RH?.>aD1@2R#^X[R--B=
:1)#QLJ\1@QdG,@J>[IYNQ_PSPDBD>Pa8@82_GSO>bCaEJ56RT+;E3fH9]T?eG_,
J\;]<\(W&0aQ1KMB^WU+:X+eC_=Q8R7bI:Q@1f[(?AA<CI[V-M>_L;e/KW,6H-RV
&X\M@IV/ZKP3_CGaO6d3K_JZ+WS1_D4BD>BeZSKa):]##-FKf>.HQXN4:R<E).Ac
8Ta<399+H;E^Tb47&0@Q?4]O]PBU:g_QTW4=U^7(U[_\GF)J9Z@GeFAf,7c.D20d
^S&9\:.WLc41@f^ZG@LQ-19Oc4+#&QZaTN:D[;X3\NfHV+TS)@(DSKfEPVcKS,7M
=(M8G6(e_<+K?AJ#SX)eFGfgO>C3;Y^8G+7G-,XW2@>)F)VB&M7e#1X4/#?.@71=
FbJ\Yf<@AAP8&\LALJ/:UZ\VR)NG5ML1V3d^9:gB-3<T&O0a/eJ^?CaW)21>#50T
+eG3aW[F#5.a&+2E>CC7/H]FK9#:e/L(?]X5/Rf05bMaIC]-3MK_Gf=PI(4eJ_<=
CNHa6XKP/X;+_S91@K.NfZQEET(a0)#d>23XHYd:&fF,BCT.+Vf[@XTdRJ2<=+P9
g=X@bf6/2[[F5OWE5W<:D5;16>c&1E<YIE=fIK>]0f6+Dd32KASU:D7#HKPE^?-B
-@[VBL<eV&g>IV-^e=LP57+PXQb4baU3GTYaZW.aBIdQc]IHG,ID_IPf_-14HK):
0.EB.VMD_HFWR(0-M;2(_6J<e7OJ7\gB8(TXR\;>7<N96J^2XX&[OJF=V\J<CGOR
9_])++JM03U9\4=S/b0^bR]7F2:AEU#8B1^H]RG;S5>?fB&\4#Nb<;R1&R4#4E26
WFC(?SBQXQZQ^VCLg#.Ff6W^a3WY]:=NJV;@<G_9M&9]b+^=OKKC;<C^DH5cgf>=
3R^+fT+SgNU[#H28L/QY<#[X6_[NQF<Z#YLQ4Gff-g268^b_SAPVM;BUc,7RA/<;
P23+5;VLB=PSMd59HKbVbEaB9Jf:S3LeXY[T.XcXgC7(=cMWKQa&>g>?9,=D&TY8
0)_AIV+M8Cc8YK3c6],-=)X24Z.aCf02UAA-.\&KNERL8(65J9RMY]75:PMTGfM\
_<F.a[6c_AIKI<AdU2dS6<.Idc\Z<(_5,MJG]44+eZY(L5f[FUf]XJ>D=6D0D6M:
9VT6O]]FDdJ4[Hc(Z495F[NVaJ_T0X_@I/[<ZCa9N_g8@?e;WXe9B(NId23H_GKe
]JgXU\M>YgZ-e.W7IM_:g>GG@]H_J9U,2C9B,9f#US;CB=MVgd__@N6C@YAKW[#^
UR9,g-BXcGN+c5Q0QJQY_#Y_[#\feZ^.C016I2/ZH^C>4C>([M_6J-0I2GPNRK<P
3S^1><>G#7G_:TB8<BTf>=fPc=fL)OUEE)7-25VEP:,0f0OL[:U>2:/c5J0I7?fb
dH^aVQ6\PIGD;@LNe19P.)fP6$
`endprotected
endmodule

module SUBMODULE_2
`protected
JgI56M=T1O9(AWg.-e&1;>UZSEAb#PCH@IaZM@N:)E8X+@9,6L)Q+)J@T;FC[D\/
\[.G@@WQXaY[87Qc/W[ONS6R],8E-<-7JO8<VIg^94^\D-aEL;b>UDVC7:0P<Na>
b<Q75N[b2,JD9EB4].F2e+^MTT9Gg/P#d-I#9#gIg84(H<;8A6.71&O)g>PVWfQ7
PJQ6OJ-1ML8V/a6NY8=I47F]7[+&OOP>fK^,F2]eKS]S:)gS7a?+g(OW#D2^HIO^
BJ+f/\JDFJ<GV[fQ@d]=.8]K\AM:g3L_^+1+M]f2dCM?1bEL;A+Gd)V&\CSE0E8]
:Ub=?>cSBded9T;(0a=DVS-..RVF=a3dY/\VJS+1F+Z<P2>,Q;-5HDeJNf<20fBM
4=I:E4f0AC-RZ/6NaYHRA;<>\^UD+SN2-8\]Ue1#)5M9VT[=/,>NDBB_,7HcC+CQ
dgH[K;4W_2CfDA52XCQ-=;/F>)>ZS)LLg0@RV/<_RA[<5d:/[V.W7+EF/,f?NR<V
]_>/3C-4HJ9_Vd-/9S5d70R])_DH<DQed&:F)^\K/^0RdfQDVU9PAFOS>PY<O1Bb
<<QAQ-=TaQH?7ZX,32MP_^-J>=+^X(W>&1C>3VdEEd[Ba7FL5FfF.O0g1\,24:@4
M9;]A?L6TRLdDPJYZR4Dg3gN1#P3[=I;G\>HTY_[ETP+3J#DfM@:Z8e(9:LgdYH6
T(5KCH/)bH<(>Z9JGMLAGPgN7$
`endprotected
endmodule