//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2025 ICLAB FALL Course
//   Lab08       : Testbench and Pattern
//   Author      : Ying-Yu (Inyi) Wang
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : v1.0
//   Note : PATTERN w/ CG (cg_en = 0)
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################



module PATTERN
`protected
K@H^<0GS60;dE7>V)=?SY9E31DUVb103Z2Z>B\C>21&?_,UHXDLK6)FZ]U[0?@,K
)7ONT08X&EY5D<;H>B@VN#[8BJP)ad\_J3/23[W-B@#0I0DaV(eQL\FABg6cV:\f
J4_#F]R(LRGZ=2(E8c<=Z4X/SgJ08Ifg(8eZOSbU47SF_^^1Q_4(=>.e+a4K5A-1
PADR<N?^Y-eFRTIDZ?B3-Q5=f1EM+-4B]#PEVf1[R<TeZW^DI>Z.Ne_&b0Z@GI\H
O:dZ_]XT[Q7/B,?^FT9@_.&S+TA?e1ZYTg-cM>)D#5?6Q)Q44NIeg14SL\e8CfZN
Ld&NdD.a-]Y3/W8HVO_DG@G[^ICIdX?8RSQW6\24.JL8J8D)8G8f#,Dc-,73FOUM
bU;9/_2BOWD<WR+>PADFI_-+I0_Z3/]3,G5_[fSVC@=6dP0Xf8[(gaaI=T0<[Q(7
.L:OG^R/>1)dTWf./LG>G8_(QZ+^10cHR/&7Ed)\@db?EeR1_ZEL405M<JSb3;WG
IMLQ:9+O(<QLK<F<fY9E2=Y/DW(7d>)f/8F7NG1-S[401<]0V]^3dNf7gS/<O)2Z
R/3O:UN],+cIL6GN.W)ZIAf2K3#_(QM\#5[]-6Z,-d#SD8SFR@b<(838aM#KD<^J
a:9-F;@H6WR[KE5XWB_N7XcLcJP)LYbGX)a2\F6L.O\d<H=efMG.F2QDG;,2ZF7I
/O26LS<D@:CO;-1]+N&;M6XA<2JN;P4JLKLS)eRC__/N:)DP/JR1#O-[@_7Z7PTd
ZGZ(2IdUXS=_SPgc^NZUK2A1R)a+a()P2O)<<1.MA7g(44Qd;=d+gd4OJb4dXCP?
@2MK=6XdFAZY#.A<,G+e-X9+-LCEB/Q;2+9+:D5+-)d]Ub96^^d\I&KKdf9-:fKX
:g&?.KFG\JeZKdQXT2D6NIAC\CM1-I\C@#a3>:;CNSFW1-6M0Fab\45A@L;QIafc
S3@+-FFAST16DX__)Kd72DX,Zf:I3>#)be[2H2,EAG#>]A,a?fcSM36]B5(/Y9)N
TEXN9bXS5,>;S0GIS<&c^PJHY5#NaW?a(F+&X?WeP33-Z<Za=\M&?__[;f_KKDG_
F4#^0,bM(QGH3GZE2GRBKcTLa=(X5b0\4E@.F^_eCT2gdRga#+5ZO?&;.I8GCg<O
.EeH1fH+c)&>@:ZU;2>g@1YW),c<8-2fgH@gS.9gHKWM6.Y+HE[:ZW/R2Y90U[IT
)8d\4Ee+@Q?N6;,=)Tc57Hd29^HV)ISDePPDeQQ.eK;f\8#?_SNd/Nd]Q0I/K8@W
^G7?^FMUFeg^T-257]#FWLNW/)bf=/1:?D6g1CD7CYFMOZ08^cS,^RI5I,eSbC#K
Y=^T8Rb-CC&;XM)ON,gLQFL)0<cLRW<^_6?/Db,J?;:;-=_BeV):V?3c(<7:<)BE
\?Q?8YP2U^M2c3+]fO1+@1U_OL/(/[/\-1)d<LQ\2Qf1Q@[5aKg,b;447O8#<8\0
+@DAS9KJE=EQ:>/,K-\02^J0:+&cU9Tg_,/T@f:&?\dg_L;HRV6ID8C\bH>Q0O>6
CB1BF17c0F-5Ya6QUVXY3;.ZRIXf_VDVe23K6&QJR^TMV.1]2MS1,Z9&Ze>/-g[D
Jd)]O<^B6QEe3cYgDB+BBC0OUa/O-e/^&bI?<H=1ONa++Y2DV8,+VSa[Z12?YO:Y
gF9X@)GEcZd(fNAOaBBRULM=7=BHOBLWfeAT3N=9b5C[J5,G7dIO2/G&KN6S>X]^
(9aKHB+,0U6K)X3ELU=E14TBGPIeY0=@2BD-68T#I?V,,>e<=VLUIZF7XTb^@=A;
eEfPD)d9\.Sc;OZ#TfMHFV=LL@-F2R_>)Zc>JLQ=FK0>)Y=g\7G&L,50F9gYdVD3
=e/YK<((0&PA<3J0S<L<eMZ8(Ec0RYDG(V=#JU)<G,f=D?VE<NSAE/RH5e>3MED<
N;V^L[HXfafM1;<..X6(Z1N_J0_]5g[O=N/=6RgaZ2Heb8Y66c]J:RIgT1+g\fT0
>N8B?TGE^V<L-S_68(U:,GLV,=?^#66::&49g?gW-IQ69SO)DL;,^05E<=8^5,D[
Re:6)/E@;YS+RQK_(fJ2K67Pc22cV27W5eLLP\H)X30C7d:,_bL1f()O9#>05I^)
c&f93f(GO\H8J>9FG+5cWbdL=5,J5I-dfg6,+E&b4B;9?B\D?;=4bb^1:DD#Be13
FGP4/3/].>MF<@?HEI85Ra<LgN[.f295cb6.<LY0V=37:a593W[a7JDV?6X#V4DV
#FZ81MAg#8b0QS9(R03TC1AdL(g+ZB4EY=TQCIF>Q:D;H#X13?,7[Ha]d@NfFELU
78g);f&P3_RD^d<>&;AO94Pc[ef?SKV<:-G<6&fQQ4ND2;IFgObT-dT#VYY>FXUb
=<@@IXeg[^Z6:3(Lg;F>JOLT-V,\KG6W5XM@)O_I7U.[.?5-)?#YRdV^J#,1e88W
:HEG/e77YL3gV:D>/:Z)#ecY<8C-T=1L0)F5=g2<=gLef>He;]Z0baJV/DHTIB^f
bPC&33S<dIdc=Y@9&\cb@J&)L^15@b<AD#+V/7XIJ_/dDH5JQ<:\B8EBEf7e=R2Q
Be>7^T-K30a(524>.LEUP=924)VX(e43JKCZRKXNV+N_3PSJ@61_GaD>_:FEEAK<
gbZfa??#00T1JQPfK+K[M40_B8P8,5K[IV--^;?]);<6BZLV7L&]H)(I;ABa@/gB
SQIULc0QHd^OeLMRPXfcS5U5RKUSA/Jc@d1D=FOd&<(44Z9eWH4.NLDRTTN;;4]e
J408,dU2M:fI+C:dA0)]_[Z&/:e,3&3:0K;_GPT#bDfH<[c2DA8,8dG0=H(H:YFB
=?\.;2BIfAATADTH]V._/1gTF6XE.NII9FFcJ\3;MCR(eMVXGQEGWSZNG:,=-W)e
]-MbIC_>Se)CT>Fa\&;9<1X8O9_AWA5a7&)LW?2D/b[2LU]#B5=#5-R?#aLY(]e1
.Z\H=AM@((0J?.eJ=JU,IL7A74KNHT9RSe(6Z3SOO86&]Z95_HBH9FJUC0(@fe&B
MYXHb;Hd4B)[D@H_)S5GYRS;ORYW6/&C<X/&g4NDdADV-M4MQ,3fbZD4f_DC&.K\
5d3/H,Q#([MZbU\?a09BZ05A56]MW21?)KdN]C>L=I84fVg_16b3JIQ)4;?..aKa
f-E:7O;a)V<AGBFDAfK5>S9;)Z,7GB;4L[\X(J/@@:5\,V]W3Uf/J>N\&]<@&,G=
X+8-(E]c3T#SC1C,Ca+8Q:7@T:ADSG.[VXb[cc&/H5<2@>:8QDb[FWU0gH@Z)]^d
Y7G7\W70202:E3_Z-&c-KISa65IMb(E9g5AP>f#F#JX+P-f_4RM2Tg.1PJFL7/&F
S-^D1c08,dH,>&gg?Dg[2\N)S#@4<4X.T(G@;bE1-/A<VO]gGV_,DVVcKe/XDKe4
-DUJ2?JedZ4KYA)fPRL;MNa@>Z-S2Z/.TT.DYJSdYX^=<S7FE-(+;&8\ag07V]@,
G#J:^MMR2)6C#SB65GU\<W2F-g,@TDA@+AD0S88\b]K\5cD616XD^Oe12.FI:@g.
SEM<5&^N1UL\+I]QQ.6EM]?W2&8g7-VR#I3>fEHc0?3UV[9/bb=JC[NdL2BMW3.4
:cW#(Z)c^L^D>G,ZIY5aXJ4BfL+-RRQcGJOD>VMJ\_X:K,g\4Y(8+AZ8#\QOH^9C
02UF9>MS-D\eS\0V8)H\@A+\Db\86gL0)\P[fCc@>\?1-(]NURW6&PWPd4[PR>ZM
CbQ_T451:[IK:L?+(SL0;(VIf\@?K;,]Z]c_]Sd51C+RTFQ/?:g+_RQWAUJbd9Ke
(<N[7Q/CR+b4N20+C^_6#7B[>(VIWK3O?-GL0&G5,89c.C@a@OP>TN>_(A(?AR@^
1<;1NbEH]#7b83WWa<2=QNK^&^@ECU1\]]eW+gTg^CH]f2M^].OL:HV[R0QMI.GR
B<C(fIHGSU^#4e]ULfV2;GbDZg_:&H)&@MA9+<:Xb[Bd=[[NO_4J=TUObe#>;>(C
<1:EL1Q+U29H.KD?O;-]DF(X,b@N[Z?J-)2<5D:D4DaLFGaBH>B676W?&Fa<X/E:
?CYd>aX\O+@1F:Z[NZ5d_d&)T/WA><?_I^+WI_QGP6a1Z>S=\+:^Q&EC0MFPce=e
T-WWbM(Jd\(5/VK#6EPSNG]7bcS8_97.OE<#@Y84DZD3/P.c<&P#9,=;8JU[#;CF
X5ePS7ge>()-=YBH86\<5KT/VL+@T>2_8U++E-7B;WMXbK1H1>TN-eL+?GHU?eH4
=LHF0E4(>66T/7]UPfE^T=]LXBEAg3c@cLXg?(,;DM^;AL/+3AIg\V;YZ;_9_V\D
3T:.,8D>M2)eBOCeJLW6-5:EQc6L@V(PLA3Z]7;Fag>WU1W,6EgT#;?#?7R\2UV]
;C=_8@4g?5C^5+&8W:N9=,9&g7XgKSLNedIA7DeGSE[<87L:-3\7PW)L2]6MLLV;
WZ2JQaU=A<=QQDKMfN1XS#;.\eVa60dcXH,XOQ4-C@(T.Pb^fB,/J&SM_HJYVAB>
edaUK^;45<)NbTT:40[(Q9H]D-:?UB0a\#cBW/=F.^2dd1-2YR(D.VZgI-/]]<G1
0LX&7-A@?Q[JK\JM//Q&IQ]04)G\BZ6OF=.>.IY+ED7Ab>=6aG4C&eG(6C7cKf;3
&B_TF8<Q5)9-(Y6K0]@8+^-a?KX]3ba=/B.C9XKdN17LX1@R=<0b;P+[0/MVS2W6
[eM\_-.MW+@]VYM)NRGSYF\_(#]XMFSNa[1)e8JeQ>0U)4W48FNFWK?UUFKc<P[0
Q=7_JL2+L^Q6?.Df(E^bOeK,]P7Q684f24@7OY;H>eIUTFd0LW>(:/fdbK_W#_d.
5b>,)-Dc;6Yg?:L07De;\b_[LJ&0I8:NT0A(g/g?K#/Cd:bU0b0AB_\4f)b#/8SG
PAE\fb+?f\75K7#/M]NNKc3FQA4&6/HRd309a2HWIYQVeVW/WRMW7T0O\P18S(T8
SBW^^[]XL;Za(/A0NU;H+K\NU(_N3:P/bFaDMW8&)d58=/:g2fb4.59Me3KLO_fb
^UeV6]]@,=-R>.#4<VRJ^88VF@HQ8EZDPF?(0F8gMdbL)/]5f+La3;K9\U5L&Q.B
2;CK]TcYE1^@2#JTC[#UCVf4JV=237GH01[3F1Rba_CAQ\+3bH</2K+27A]?BXdb
@.f/9IHKNg8aU5+&ZAUOIM+FT;_a-XT-85_H>F:Q+LWc?1/R;5_Y69HdA)Re)^]I
F^d3,,D;:1RD,WX54UfIF113>@Q1W67)a_\bgFSUYWE?@\0<.9,2?Ka5-C&a@P;G
gY5g>5)JA5>dc7;).;W2Ze_X_#R;@#;JF#WU3X&8GY@B:c)[b>LJ5gQ6f?S[ZN=^
b,8__][I.YL6e0BI/6fL]P-]<\.Z?Kfd-WT;[U,_U.U1OUJ>+,PRVW>H#dLK;WMD
?.8],WE2cf_+Jb7;LUU0,,Tf+)H??I;g.Pg):gG<RKV5gg;[aZUB1W4,=4_UE=fX
,bN5_7MWJ^VJ^)eCA8\A/H/2Dc0\H(K2&GJ0IKI?3-c(JRL.F7TG^a]5U.=<c-eQ
(50c^,[<ec&KJb#Y9gBcP=-\Z]9Ke#O0#DcLVd9Ab1H8&]9\1;2)cP:Y+,#7c;9\
?+\AP_03c67_V7KC.N7CD;HB,)WTN8H1YJcbgNWe5()@DCHVL]Hc)PaK--M_KRb3
X]<B@@D/1U8N0dAVHbG@,OYg?G)?(+[7#./0<54@B8IB^Q0]UE)EMaLJ0)USS@e4
VBR2gM>,\dJN[D+/>#QU\\L+Y3+f.gG41QQYO^,-MY.&b=X=@0R[RNY4Ed]NTVc5
3IESccN/-4-T)bc95_8=ZU2SL1,F\E5JT^cZJIO]O)>?IVO7RSR#]^a-\MQSc5TN
3(3/6;)9=9T#;8Mc<BK?XED]aPC(+_0/_C?0)[&+/7R@#H;:-T@_=E.,L=d<F-M9
\_PPO7Fd0Fc8b&,?LWI7NKZa>UNKEMdFPf&OFaQ8>XB,97)G-AbZ[KR_V1CXXUTP
e#L11[O)VCW65D+-XLVGFG3X:REDM)EBLAYFWJa7MKJUI:EMH(SV1cZ4\;KZ/@=A
EB[BOZ<G_U)JKg)_1X+=S#8X&V&[eXEB[c4bHQ6>:+OC^<[O?SDS1EK9g2@S5+BG
?T1_><+I+J6L\Of_eA?&>9KMTB_>Ae2[)Z.]0R0OKAOIf,^KEJR^0VH1^<].L#\6
=3fY1A4GV]8X[[a+U0H)0>VP,aCFY1+1)TM2+Z_A6)UAHgPTZ4XAJ;G=NCggNSVS
S6^,>&#-NcU,Q?6EE#K;?FH=8_-a6ES3NSUd[MF7+b9/@8Y=a7-X[M>.;/QZcQCA
[?RNZ7YB/.:fPFfD+)8<)J7FRb4^VOTafdW=I5=MgC:LL&U-)/)g2UA),F.)]NKb
V>aG,WG#eTC:9(b08=bK+bE4KS+&FfE\GNTV2;P=WL8C1U2^HNK)(e:cK+2@OR_G
)6<8390)5O4)b6H<fHJTQf,);LUP,:ZK-9T8_g/EO.K4\__8>4</8_XIaaf^K#X(
BFgI1N=FGOD:aFSI5L3FB(R@_^BVN?>EV:(&a<[Ia3Y5PK(FbX?P@01+/Q^A-aXJ
+Nc)\&DJD.:Q/62]Dg)5M]VXW7DJBA@RIUU;[4KXb1ELIYZBa_S4Y1FEd(eSgDT/
V34DPKU\M_I<\EL-I6HH#A70GO>(a:8M/,DZT0R-X_1W#]0e]R7K6dN\b^W8a1IM
6RZ&Td+<?_(@AN&QccXd_&<49#Y:&:H.+M^E+YJ[>P2W)<<05Y,cKV@IeKEd7\4?
L=#P#K,]>ZHJd1+7Je4E(5RHH6S,,Sd^]c_LQENec[QSM.]5cga-</,FDNJ/8W&D
\:OR-.L[abN?VaL&Tg4PCd7PDJ)b33DX&X5M20d__Kg0ec[;@U946;9J5B9TXfT>
I[f7N;S.4(_:@e,]059Y&TU\N7Z3G#;0LM?2CR3W4gMRWS-b2W&gg48>H^d[RBf+
=)NCM]).8\P.a8KN(,TK68dTY6&.>K@AU[?#a0[S1-KQd7RP<^W2JR<RX<:Vd69.
K,/&(0PC:TI300NK]8AA[1,I;=7Cg0P9-F=,^IC0-3/5b:N1C+\P?LY;58GGS+c3
.FYCg5@CdV04cP.,;BJ-^=a^T;MggS,0C#/MSI4PXcb>([9ITX>?&#L663^\Fcfb
ZW7J#a.3b8SGb6g12fO4Df<6f)c@Y7929Rf:AR^BgcXN7d^<@&:V<Y:C4FL/YA;N
\AI;VIA8UKP:dAERHKJ4YDG4=BIUU.N4_4b[I,#Fc12_a:.FKRLT_^V:dgUG6I#W
SI4/+VVVT/^G>a0E]/B7A9.0:PF1=\6VQ(SAWe4ADW6PA;I&<c3dH-LQ;gN6,M\C
.5=^RMF=>S;4DPQV#ZUaU+0GN8_O\54dd<=[#Z)0eR5-]E;adITOVR:[J131+T[9
NPS-BERPcA4+1/(Ib\:,Cb8dJ<+<)X)VLF=LTMP>BCfWMGWO08O/XC.Kd@)G.63b
1f[-O<?RJcX]#=4N.;VcY>dJXHSNBM.IF/Vd2OZ_H8??>WBfIG;SL-_WVL/??.)G
.&65.7G_S?,4EVPP<GW&E5MP4U3PTJ@7#(E+-1_M=\63(f4\=EeD-ZQ\\?X[W(T:
Q4_O>\OG.O7NF-<4YdE,P@B=P2cQ+JC2c78XG0cCQ32>RaN^28?f7YO1)YK:D:/_
SY7aK6b-T)5U(M4#CTZ<ID@c/H?FQO^W3cC>;ZTF#d0beJTM4_UDP@A0.OH[;deV
O:S<T?+B.J2Kd_\3_YW+6=NPQd0,fdb:V5EfT]]dPS_K6FL#6I2X&?e>G(V9e)0W
?3RVeMB.cOE5H;+O7aW;5#\eWEIQ/?KbSZg[3VP<OSCCYEIZ/Y94/IT?gC9L:NZW
<&UJHM<5a8L6S=6@@GL)2KK\B]+fPecC59bBL&]#Oe7cWKga7YaE7_D)72Ybg6S1
W8@()WJDL.UgX2[Q(BY0GC)5RF[]Dc_MSR0dW^QAUe,-a4[B/._\E_7N9@)I9^KW
:Y^K&1JTM3T9RB-L^X8/Mf?.-)938E.5N([NGRaB^a<C](-)Dg,CNeC.0GCY_=a[
+L=U_d+C3BQCJ+a0OVC+MdLZ0=-3Re:#,NTSX>ER?H.BF[I[69^d^QG]G_+edN4?
ZP.5\Y7W#S+W#<^GS#PB]V9-B>ZZ/G+1>K.:G05@/;dKLSQd@Y1Y0U9QA#:AZ@M_
G[)P;5e2MdD5O;NV>G>d(Z/a5K=:KIeL?XP;CQLFGKW5^93Tg)bC\JLVZ8]DID>f
[9Jf[J]RU/VK&N96fAM33+V_WSefaKaCP#8.IO10XX+<>=cUIP2#SCOM2N3f+?,6
V&bCf#+M\dB0/bLe-1eXHBdf;_\6=cF_Ic.;5S7H-JN34T^a3PH\OKe/H:W[[,I_
D6:]PF=IE;JHE.WT@,EbRNMC:6?E\BaNN:Ne2&\W?2>LE/EPM24H6.4L@[+04F@e
)R<cUQ)gEVgQcFYQ96b,HbY9X<UFBD+Y9c1.N\4W&W12dQeFAcdNXTN)YcM+?AXd
MRcM.ZA=cW3TATRJee/3EN\AP2S,dcCRY#4T>(b7QGY1P27AE9MB;897&HSOD7T7
^92C?FAJX_aPf(ZUKbK:+FI19X:HF&0;1BS5/C\M<3Q#E6Y\9]O<X4:?aS+dFcX8
f-Q<-,2FP=^,a[52\(bSX[H/6//WA(f;?dQP1WbM37e6<RN-2W1#-OL&I+^^CH\R
CcQX[g.:MG9Q)3QB(<A90=7A)P58bXJ8&9Cb>?UWd>KK;3B.Z7Z?;Q)Z5,4+H<GU
@.9ANX;;K?@@4@A(aQ^fJD//NCb,JN6#g3[[b2T>H5N)1FK^TR7>]S)A7[dM-_R0
J9:Y?#^6e<(MDWQSO/V5DKBPdg[^7KXY+[OL82<R^KX@<\Fc9>VBV3a6E4g;]:\f
VH@[+L:6FUPXS?#R;IdS9.2edTENMRe,:;Q)_4=Z0)4IRgZfR2bF+^MgaC]C>X55
<6?@#cO4>1@7B0-88e@e97\_=4T@fYVW^84cZ+D-O1bE&dgS&MR>RQ41^-X70YfH
H&G>E-.(=5fJB]H=-\Y4TX5AeFd6&FdB?_eP4XGDM\>Tf)4,M)A_.Rb\LHTKC7=g
X)bB5;>\>@Y4_D/7VXNXfP5>SD7a0&8cO]^gX;IM(g:M&O<g[>ZZ#,bdYQ9@LNEN
^#-FGbV+Z<]d1VJ<24C>9X8A0PW\Nd]GCY4ZO@I>FQXOR81RU0W//,Q.AH-H.L,/
.+RU[5.2;K<MT-0=/f.+=eJ0fMEb,>]2_dL^#(YPHUK..&N]H-YS-]NH[Ig0G/<_
GY.9];^(:AY#Zee3eXFSOb[9O4DeIO;#A(Gg)^QFSY6/KcZH1(dXLI[+dE>RUBNU
#3J,N7/c667:e2[3-4GGMQ46JCG3SC^g(J,RgFQd[HRbY^GM\<9HX8W@^1H_WEN+
4/LYbSR=[:DZ3+)F6R89(0B@C#\:/7LWcH#(N?MS#aC^.^OS,UWS_/--bJg@2R2H
T\D3N3A.(C8.N+aSD&)K4L+ac=NcY<Yg)(9fBR#L(d+OMeHH9;9/>J;@)A@WQ+8Z
=fI)1&2dIEE<fS3[6E]1C6P]=YAG\gdV?c&RE+ZG_P@XWUR/9@?6_<P2+g:a_U_>
Leb1[_=3+-Y^?M#5KU78&VO<Z-GIGS?.aNR7:2\c;8O6-/->Db-bO7ODO@UBPZ05
JRW4A[g-65a#D>gBCVL7C_YJg<0IMWA?@6eJ4aeUOZ-&-@JB#f4DY/[#DNO&T<(b
,6c+V4:)->L;d]U\,eS-e>8(UB<9G\a?F1P>?/#+f66gI5I,#fB-2=\0+dRgL[YF
;\OF@ag]MDLP3Q;FAAO5cdNH66/Y+/1CN:75Y2,dAV-=I,9?U+YO1)a>(RU28g/,
_S2:]5b+XQ5VB5LW;@I5\3NKV.A@KGMJY^(YUaLW-PG05e036gPGKf[:G[F_C]D9
^][@N;5b0);:K9)H<d\J+OD@,g35I[)7=4)ZDP2,PcF(L9W8W4bR>;MZ^1RKc:bQ
/e#T5Q:^[WA-#)>:Tf?46:BE9g/U-P?_4>BMC7O-e2IN.F(PQ\;SXMF=7EFJ-;g>
TRb99L5E&D^VbGV?TB.eY&BYIIMX@a>>T(S[>W,+c_=\ZAEN^bdCcA5]MRK;6R=A
RJSWe7F6Z2a:e_c:L929BK9b?aZC2HXQ;O27SH?F64ZO9S-_.aUAA4_T0Fc6a\U1
8;5cR.J#>71S1YYKO,,7:E.#M0gIa0E-T#ANCYEXTLWYQCW):7?C;eT+G,_QR;N[
Ab)LeMe=8;BER:&8cbJUO&S]79fd1KY8SA#NAMN^eN4[X8V>.d?RO^OJVeS5,?(\
gN2F2Gd.c]_U\Y7@WUW0ILFfD-(@3ZN:6RMcPb-ZJge-;Td^GLbGW9B-OKJ1W0FL
WD9DN0-&C,\]NU=bF&=f^cLeCL7-RN(#<^Ve\D<]\FH92Q^T/B)1e.KOH5N>L[(b
56,P+=@60&f?L9Q\7b7;BaC?:A#NKeQcDK]EEJ,<8Z.3<)1W=,.e^3@#XP.J-<D&
@)5618CR[YW5V6ONLD0AGVgXgG?.0748W+KB&ccB.@6AXd==SEMBF,L1Jb#VMD9,
3bXA,B[f.,dPDR5:5>\[)e=+^.IK)BEcb<gBU]VQD2LT20X^76/1?_++56#bM0D7
5>cXgUH5#]b1d@a_)a[FIJd77DeWO--X5IB/@Mb)V(]MTE4IV?70#\G^YOMHE5#:
SFLa8I@OHI-L&1:VdcNQgG:fIT#71B>T@1U)TLZ7bQIcf6R#CDIFP&&P9bS@PS<S
&I\Y(;,GcGGG2aDa-Y(:1SfZZD0=M[f:=4S10MW](+-CMCVE<RfgFZ,X728Tc8cQ
.4C8cWgbNG(6AC@.CP8.L6X]g#0P2#K]K?65faYMQJF0c;QK_J/1:WJ])CB9ZC0R
WQBLeR^P>L4LaJ]]O[D#5=8JGa_-;#a=I=#H>>WOD2FL/_f#@TR@Y1/gA)?421D_
Y5@M?K=,bVDBZSL2JRAX=aJYW)_YOeQ;,U1ZGQQ?P4[1SVF-@0WD+9H?ZeD=MD.D
ZOb#IDIXaS;7IFXB5g3S;B#dd[Lf)95?:YPeWTOBSbWQ[>g(@Q>7VI8>A9X6dPVg
9[3]/D<AMB5FXVSNdf;>S4FfMZ2<=L,GW@6G5FaQGdCO.9C6O+^Q]?TZXSL@&7bZ
21#ZUDB;KV;_8J0M-0[\WO,^faR]HBcL9@I\75=#3)/:6#^NbU.N:>FT3OBeZ.OP
dG2D@=F1A1-@TW?[59BR)NNJg]?N]^V>33=@)NPKO.\<gWCBS@b=HOREJ-J2WVXa
)#ZHLIA6d[<&5MSAW-J75A9=>,JMY>LY?,WE?HHI=Re4#de11#Zd)bTS1JH<b>2Y
ab8KL7P[f),=Q9bC].6HN&,L3bEE&&Dbg6eA#6)R@.<b?@CS0L2[D&d2Z?@g\fe8
6#1e_(cG^;#C5&_DS:B2L?][J.09@GI2;E2>Y/cbd-0-TV-64WDNYHWQYF+8_^5,
A<@b5c(1/PJ679MBg@&FXdQQIAaVILQLB&;<5^;aN-cWc:]C=V4F)JHWbR#Q7<E-
/G=AUGQdAUU^;DD8W]NFVR=d41K==UdMNX0,b9((5;(13b.D/Y]c3(J>^AI7I)@?
C7@5<#&?c-U,LQXD64&1>+=U7XB,0S<<XL-/bN<9F^g?##-Q=Vda<;WENg-Hd?@]
QXPZ_V9UFE[gMg;FK@@(1:GR)Td]29;fU@T/W/bOP/Z#8.Ze44-AZMb\<E8[bUbG
5ebTDAF<5DgJgd@/XQdA(Z@2[NT0?Hfa;f,IAg\=U9_X;#G)X;))HE;DXcQLDJTc
KKa/B+.\dMLcRJ=_._;1N(;&.7CT?+9^AARQeQgNCA3D[<gC<;;;_\,WUR>2Bf^a
2VZ.f\8SCTWSM92FL/.S6Sa\8L2-_FLBTYEN<(O2@D??QdN1,.8(,1_Z=MQF0YI?
U/:.1&8H>J=G\gZ3ZC;#bc_1>36_[.2(=CccODI9X-Ug44-5N-:aIZ])_])@:0O\
NJaaAVR]UO4#XQ5X:(MM>S[[:@TU8)aD+eRJX&#DPJHJ;Y6Oe<Y<c8;7_5DeZWS\
d[Ac..b<3U\)8[=).^CJAT-1MO[<\c(LCGfe9Q6MfWcO21^;B47#gLf64_X8._Td
-3743C+UH+(-?HNbc1#B-?O4C(f83?aH,76AZZ:[I0R:JCV3#M.1a0_DA4^YWP3c
D.QR#JP/[e&Q4O:V^FSEA/P-#Q^\R/DBKGKT,RWV1^ce?NMf5?(5<5)6^HeO;8/g
=[g?2JTAHG:W,a+,R/Y(eT>.0?J>.^8G+3V7.^=NLaK434^KTV@#G>W8,>HBWG.R
K:6Hb\:9)PZ8KWS76Lc9-SRYMd^>P.HU3dBFA=MH?7FNC8a+?B:.:</<[Y/cT0)a
TWSW/I-S.:G#Jg3(b?=bI,).RK)\bP-6T]H(,d@OO[AO27bVWUX>Fd:d;6)WbN^W
]OX)cT3G<.7:)BK/VZ,)DgFSbYbd>/X\:4E0,c+,](HH[7^+;WVeBIcB,#+H3[eK
O87CQY1<J;bfBbdb(OB6+BcZEK?OZRcJ-P_V^HXR<P<]?/&Z^2[T3[E;1feaBDdb
IZ#MD_Q?VQAO)O>V6BY+?=<aNg/VSfX^L1+WM^5MS4?^c3Q:X#W?F(K.,#e6Ya_2
:F&+7G@gNBZ)e>1<=WEJa,0O\aBN8;G[S8CWL=855Q2_\_&FKNM<:ND,V[ePFK6L
C3d;IC9F@3E624R66:RO<BVT[<\2X^]<+g_fBJD5^(CQ5RL23P<K1SMH1GG-8^@@
#82@d6C2G7N#^#Df7aU/?:cOG1,GJMK4S8C;=<H8dGQ#VL9g3b:PeCaYD)a2cSfX
I-b[HYJ97P-P&@AEMc6a:&KaC2O]YQNTBd[VRdKZ=:SSEBHb::T.B?)OFX5YSJ+g
4H]Ya2/a(P_)]:U_.bNBbb8(ZZ>)aQEV6e;<L.^898DN0KTfZ6GU6F;W2/0:Aeag
e)R>F_U^QS(I?=Te9HW:8g(WIe26[9^@FbBH7X0E6=.#,eVG@,G;g[TNgF[_c8dL
23ea>TJQWOcSDX@\e9\C53+c4f96.;8\>c&67MW/:+CcJ=)DfMeVULU:X3QY.YeY
6MQgKUU-)+E^fgO&UE+KSA?G\Q:H)CCIPW\PCgdND9CTX9X)1@=_W,Ue@f>-U/Sc
YCF+U(6VSbPW[(T,Yg-HVg(4\H+b=&Q>0+B[;W>&_Q]L-\:CSUD8b+([g1S_10g9
(T6;<<S0d6:g58@F;R.X\:-c7MN.2;Q[WBWL52e-aAX-d3U;E0Ia+;1=BX3WPfL6
JQ;[dS;-RG72RRcdCb,N&,>g=TO(9S8D]U4Mf=Ua+IUQUS:ZBB^V[-?B-4?e9-\)
8:+b;LC>1bd,f/dVHRP2.<+\g9]3DDZ/C0P41Wc7;BV8NW20QN/d/#_+BIDN2J^.
PXBXL)8P+a3<\N60D?Qfd;[ACQ-_A@gedCF5cY@,MZF;4#b>8Q^U;3OFT^;AC4A)
-VL?=5>9-Z=H.@?-94/\-dV/4YVbL3I8C9RY&1_efV<Od=\:BLAPS^F/_#=YM>K[
#fgPTNfb>L1J?GB_IOHF-_3/eP+L]0A#&9_7:G8JG7KHg(3dcX@XW[\EUg0:.DGF
0&(V#=bL6T;-(W=AX(G=Q6cc83+VG30-ZYJU=\caAfVH^LEO4C;TT.U[J39S-S>6
D2L,;I_9M&FcRd11:.SD<([/YfTa0F-])9H9dSW=Ka0(?R<1O8<&1>8.ME2\GcaA
/bAeCcRHV&?_;A+;J#bD0C)_DA;Paa,CcSBT#GaXK6KSN]0RG@g=]b);DN@d_F(f
X8D0.<@bMWYI_(Zf@JG>a#B5JN_[(J5A^YTW/JB_b>A>8U,dfV,e9c>#&-2CDY9f
C(^>2aUR^OXLbJC2Ub03V6/)&=E@O8RgND/Mc=#CdAK9-e9eZ#PQC;&0EVH-W01)
Eg(GJTE0H^I_N0+f,W.\OB3T1;9da()_Q5OX/-gZ3ddEWOXW=E,(<B4:XHQ)\]U<
IKX)(:FbW@c5cN6J<\2Y)XVMWXTN=YISTPZccQGa(>c@31L2d5FM4<X[5\\B)O@D
=&fG7N,<]U:8MP;bN#C,cZQ6/1(D8<[d#(FVC<V,7H+Z]NKbTDR;S;d];/fcJf6B
&3AYNCH#b-@<VG3c:-&gJ);,afRRX9I/>4:^.@1.KG;GG>V<cTW3I0=WDFA#^=4d
HU?gJf,KS]eC2#@B>]H9Qg8<ZcMJE>e6;L[fIc4/EDNdH6cP=H]598U58-T:@C5O
J057c^Vcc5N4:d03gA(e1Z0+6Z2OAC&SZ?#D)5E#:_:OZ^:7QORN0F3&\[9S]91O
R&R:G8Ye>U8XFg3GQZG;GAJ>BV5]e_?&T>f^8<C[VT3T?6MfGOPP>S\=,=bH15Nd
3(K?#/A]I>L=F94X5ROVEBJC1X&PF\\^U3JTGK\fV=M/MJO;P[.Qd1Pb4W]1/E@P
M5_3-2+KDeOJS9L&M=6RM8^eGQYdHSH6KQI[V)(MgCY3P?MO22Ge[L-QK4cdOG67
BXLaR&<F:eN5;U3/?XAedFIO27D17(BZ?(Y0&XY6g-RC,<I2A=2N:H7O2Q_Z6OXd
U1aWb>c?]b2g_9dbZeWPM0Y^A)ADOd^CbOD0f;BWB?.cP7De^8dNaYg88W9^UL(&
/a-2[d=RM5]IZB+aCL(&GTd8c9A@K8O;FS\3W_H8ea=Z1?/MG@V5D61N2#;VU3UR
^]Q=L>##GRO.[b&dMJeC[]c2N[&CS_dE1^IGQFM&2F+4U=QcGGJbC462ZX7b_)QK
+?PCfM@H7U9VA._#+PEP@,<2,DcY68/f<TVQ>)\N[#1gCT;DWI\T129;aU+cPZ5R
81O4@g>#:+TD]+KfBZ7&0DW\c=>D?7I]QB^d&C46>_/E7EQ6/<dGSF2BMAgL/5N>
,?H8R.SPD1.WN78/K>E6MB\Y4\LFZ04_3fNZ3^f+<E>L37V\Z0a7LLS&ReW=XV]e
3E]0<4_H;V1UMOfPEVU\\JY7WS81cF_?6EI9aJMM;7?QU)f_D7aYRM);J1=RW],G
B);#HL:Xd4RIe-aGVc?;1Z7^#98];f+2F;,M<;EP7R.KCA9VC8-EDN?aZf[g2JJG
_E[aSaC/4P;[bEgBQFL(BV/gPN1Xa4=6(2Q[/=e/_LTgI<9FG;e&?9E]3&\9He9)
=[UA-TPM\f0+?.RKG23bbM(J]Q4SJ\W026A@89e,=#1/\MAKYA&38.2S4d1WAQ9Q
2;:/G:[?K_3G@Z1d5=E:G1YK/Q2S.CV#6.:BG&c^MR57VA-gf-9:B?P<PFg^DR(I
?&4Ng;GS5J6(]3M=X&=eZEZ[-\d8XXAXJ.5.5fcG;98CN^f_Mb_RV;+4=Nfd&T[@
-4b3QI#f)N4T7I]K6G1YeaYReEbH)J2bCK)C^XOATK.\RZW3QVP^+&6X-H35@gM(
0.b5=3/UFD[8gSS,/XeSa[DXBJ\22V3LaDI=)OcH\-M.7fJbFWY6Z9<(VX<O-Fa3
:2bKee^S/T.8D496<R8PX&HbR2J2O16T)/#G0NbZKMWeHJ,SDMPJ<f1,3c[==H-B
X(fUJO2#74c=feB(eZDC?#XK@D=K@fEI.7[;Mf]OfU1IeQQ;<-(,HB0LYKE#?FOJ
&-g.&MA7?Rg,P19K?D]NP?_F_3&:O^>9_0EgSU1VY,7S&23[.YcWNFBSPJe80[6A
&.(=/BG38M>>\DT>F/F+gJ/<V.AU_)Y;2cXJRZUPZ0FK:@Yc^H@0A0S\K]@\bbG0
D/?C5fUJ#Z.1OeSQGOdU<LNXV6W1<D_(&J,aSY>^1c<cPMFZ5d<ZK6OPP8^?K6EP
4ZD]/dFA&V6SY;9e07cK_->ADBeMfQ/_UA^e&NFg<#(g+F[=7]4eN4bJ]_[(B2[1
:BXLL&PYQB7U.M)ggT3W8/J?#C6@<;THV37DL\a-gTH0GM@>#g.QE1b;@R-:PJdW
5aPdY21YHIS)Q&YY;856K0,bPG8+@POUJI2\\SX>-YccAPWC5QfG@L6UV.Ib7A+M
3BVW[UWP:H5<fL_?IDWd,<eBR<&2.>0EgJ@;JS=9ME<S2g(8R2=A4)O-NW=^g^HH
JOPVP@eISUNHMV@V.F+?-3<E<S>=PKU[MF2KfJ:d,W<P?2DYa-/9P&ZDXUJ<PagD
aVUV&3<2.MbN\&O9CMDaCZ4N^:e/ZdAL;c,-=IBWE?4cd?>__b3g=S+1TdNDg8g3
LHSeL2F0bJL@[c#IW7)aR-dUGI;X7LIC^g5=eST/ME\_2=UX>D?L>H^2aQ/X3(;5
;Z\4^SJe\DB&/\WO+>S[MK(CNUT]:NC&D<700X^e^T-;)cRCec88,ALgPIP8&AZ=
VfLSdFEe(E9:1c,BRD,e<&.ZK^A+K.,_d.[Z[47^ICGI3WVc]g3O9_=45A)4958\
LIC\b.)#;CU^WNP?bO#ef=Jdd0(6Q39ec#SW^S#d<M.WKP4RSG)CZK[(ZO?IGPVV
I.^VGFZ^I</\5P]&Lfd&b+96)V=_2AaeJ.9aggHEH0+@<W6^V((WFQ0X-UY06ccF
/=7U96NKgAP[E:.dE0WJ\(Y-QV31L4TOCf=\c3cE=bIS40Z./,#&8#>f6f1bb,c\
&\V<ZVODF(S1?29,KFIL5MY.-0Ga5EbU8D</cI<#f]8)6/2Re5Uc/PbBLR\Xbda?
+3QYT]c1DRZ_VVQCAMbVAAMDA64P<R@E?dFHA\VY.5.4I4PU1V>;XARM&;14W#>8
2&B6.P1Q:E^CUX).;dF3\ZdV2S85RG3@N<YYRa+3HO+3cTH-AW<(CCMU89L4JYB8
OPAC0DN-J=T>D-P;_g+[MTgR7aXZ^dC0MfEc9TF5QWD2LI)IF]B2>(@KVNfgWW@\
GNQbHg]Qbc+5=T@E=.T2(^5Ka8P#I7@aO8DK3W]O5C.g>Wa3/AFZ[JaBXHQWVQL?
/<LF:/(gA^bX/RV3+4<1K+)NL)eMOPcBY23L]ge[SES_#.d#I#:g?9Bb0RLVZ5NL
TcbL.\e]^fUF2XCNSWUG:AQ;L^DMY^9AQZ5C(D3&P0\&WLGfZ7JNNW1L:48SC5MD
G8AJeR\F4I=C_DV2fCYN;:gI9(.I;f[3R/[5Vde#5+Y[8UH6:YTMTFNI2+GSW/6c
=/MX>K#B/Xe\1\fD1+;+B@M?/CHSBWYf4SEN.R-[90]]_g&9?F=R+LXaTJ_WU;&Q
Q+2_]#F+[+W/UU:B59?C;MF-P7.b\AOYf-@cY.[C-YIWDU3WZ.R/,Y.[<R1YK+^;
BUS=eC,fI:]Rcd5=T>9F4M4@]+e0@GOY6M<B_/E[P6A-+&c\IQ),FP^BHTcI>>2T
=CECZMA/Q0^2B+SYO.D)XQSOdSceD_,cc7&>@[4N<Ya#dE,6S2AA39N#ES&-U]WK
7_.2_K[A?=L&/W<4JI6H06I4M]O/2Q@aA82YdP.FVdI5J0RNW)MY/DKB2dIf^?]3
F-aK9RX0(JOW-=-fO=>f6-ggQEQg=0>YG,LJ8-I;:9D&<W;.eY\J,9cJ=.dHD1R?
a&>ATPL-a5,BX9cg0^1Z]HgLc=5DW0-9a\;+24X(BI:XC@86c@\[\1;A;HLP+JJ?
<-;[;:XJ/O;BB1+EP/&MBL=#.Q@L&Z?.EW@.NEOMU]F4-L2<aG)FD1J=@Ib5/dH@
Bb?9e?\fZA9L_^78X\7:/ECVJWVSH.)F-HdPg.?_1_^C:gQ_9JM@He5Bf<Y,4.Y(
+54)aE8g\#-\@1PM--AJX[G1B;P621\+KY@S<S0(AZ/6YO@e[PP@Y.M/5_&093WC
/:+RFE,@Nb936O__+Me__R7\IONLNL)F6>FebUc?5+V>2dWBZPALdd+Y=WX<f_E3
fPJ78f/H#C4X7BE51XRB^<da+Q-&dJ6/JR<[:,dJ[G9/9RNU:)O6H97AME2N1Zb_
&-cedWQ],:O;K4UK0-UfI&9C?KK_UA7?(AT6FB=H1dVMYC&b8N@c,4b25gY5bgRX
c.KZQRFBFIU:L=FReI#16d>2(bVKXA79aE(^)VOTDaHe?Db?FD2_Sg^PV6g6XYbI
Eb/aJ&Z];:[b;0>LQGT;45;H+>8BROSO4dVN^OUdQ][2_FOa5EEYaaSLM9VPALV/
&/X>UU3L/C+R[CY9]R#5@U@LEe\E>3Q\LZ:25R-S9)]T1R,9H.5RIe[D=1O7cb^7
CAZ(e-EbC4dJM1.dNa\#+NS2ccdJb[bb+a3STAND1Q=U+6b2R^;:dJ1Zf2c7c8[Y
OKa9V4NB=Q1c6dQTONTS=RZ?T0CQW_,KJWcfQVKb]>:Y9GXW+U7A:Ve8CA=bYE05
>F-=V[6X^F,52X]FJe-Cb;6QW[S8J5(TVaV[1CILPA<0?JSegNZRefT\R&C--36G
L9Z81(PSW[G?WGC,16OOY?_S);(WWgLdfA)@a^dP3Y(K3Y4DDeA62H3^RN\,_E(,
Hb\[L-J,/__.gI+WBRb5ZEUe^H21IQ(FR3f^@O<aF3GcYfP9T0\UY<]<_\GbS90T
_D@V;>B=>50[>^WGS(0U74IJa68?+3Q\Q.b:fW/=2bER\=2Ua6b&54TT7H,Y0[>b
8[T6Uf(<RWdgZR?VWIV09W(a+=JJC[<Kf=:DUVS?LR:H]N&Oe_]<a1SYD?\PR#1O
+(4ZH7OEQS^9[0R]PQ)b0S7cYSH@0E:V7?FIXLGY5[0eV0gQ+,8CeJ/^.WgD?EG]
EDKYUcSL66R4;PAA)aY7eg0N^aTg#dKB83V>#^X0eB9B-AZ]]:SFZ8GOV^LL-46d
I\:@1#.KeQg\J>G>[UW5R=+I4J&0AHc,21>1,(4<DXOX#A=TRDWTN03aYJ8M#UfN
^_OZVGcd3?X#FGH:Y=@_=Kc,+gYf5,Ud4EJZ30f.?047CQQXC7M<#f:+OU2B#g3M
=_ecFc^UP^IPC7Ea5XY]?M0+H=eD-aG-0&]QQDOb8g-B1W0<b(9e1bODI88J<3<#
E_4CSgagDU3^RBG1e@.U&f2<?I7Z#[c\d;PdO<51EN.1b\<<H^1JM+-SVd<g,@0X
4,9,3(@@/Y,7\#BXd&]Wg)A;K.(=Xg[W6Vb?a=1X-Z6H#[I#<<H4L4Z)CBVN@c]#
LU\3N,2@V8cg<U60+,Y_^=)U8+SCSW/F\;e\:]_<A5D8ASRNLEgW<a/O7;IJS&WK
KJMDI1X4<2,>OD06gKXbPY\2DCP=>;2V^C<J9NNL(ZJJ7Y5e^YTI;D\SFRB(cCN]
M:bDGbS]MD(<aUX-0I#2R<[5POQUJg^53A^0Z(V36\Gc<08@)T7KKN<6BEg8&)1X
b[(d,&.bB,fe2,ScH=[TF3=3R,18J#2(cbO;1^aS[\WEdNR7PA,Y+8,PK=GH><83
c8V#ON+Q3:;=(R(<A7gBZ@Kdb><MC.GV-<e2b]<g,0C6=f+3L(RZ^&23?,ObUL[T
PPZE_#I=4cUC/=BC5+@:JbNRNH6P0SLA7J2feEWQ:\WeB3N=\AH@F.EM0^SY5-6L
?6AQ#AOcWS4_T;5LY(:B:SF[K)6)DX#aSH&-TfLeB//()b7UfIb-XKXUf7N<<:fg
2<WX?dD1^T^D]/SG.?[GEOd>8[B@WQCgZW1/.A(88/E-fVSH3WLWEN\C(&<[^d8d
@CD>[2a-#,BC&dNBD:RLX\+X<)2AM;OABF7:G:K_EUPSR6G;QIK6<H8IQ:g5J#3Q
3J2__DRKbM=;_P&e,UT_<3^<Y58c^3V;I]D)cH?g3H39>f@]E0P90OH^3F+Xc\IJ
FU5-CHP(aeAF2?C+8J1R3.af>6b2gSPTb_ISeaUDL38gQB;A]d,2aZ6cag9F\;V:
ba0ERQK]b:._/+\QN^5[V+-#L@>65VXO.ARgEH0]]J9F6/#A8/E_MUdKaNT0H6aN
3026\#Y-W<C)Xc4YHL&f/[O,XUF/&b?_Q?[e9&f:=-]cb7,Fa5[#SYb+Ne(TI\M=
@dQcRAUW&]A#),dB8/bB4d\)W?_?H:_/ed\S(&-/ed6O72@IQSP-JH(CP67cRKR@
&:>[LEO8LgUg-Ib5<MDc1^6F,<0a85C/@R5W0+@c>9W);MU8,>&40=6^8QNA41Y?
AJ[D<A2ZfKgK>2,8/aYdN2HMHd\?.AILHc2^Ta,FLT\^&?QTS,fO<5\OGW&QG,-&
(5b+-S)c<NY3cBMD2KKL=H,4b,-;fIG_JDcU[74H0PAe89@?9\8YZUHM4OG:O:-?
C-@U^,c&FSNF1DAE>2D0e_>TK=M+-P)&FA231;DDUM0<;NZP&TB+F4Z]O]_g@gH/
cO@\8:^)afX:?;UD9I.TZB3_;0gH?ZWfYKM^0e)=6TT9<50[f&^c;1YJAGL=-Z;E
@#ge<cGH390L9LA^X7J=]Rd57c)<KQDFVZG15d@(EG>e_H2<=GO4>U6B6gbQO&H2
.Q>EXMS_GeV.[b+&<f&K)3J:&1J+A;ILD.^V/B<d:4O5A^S:Z&I2FS>B)f@M8N]Y
TI+7[L(8ZU_UF)>#H,YUVdME]?a3W5]O5OdF/J:.F)I:@5\_X]S7&-fY>UJK.9Z]
V8<<eGXL4:S5+.,5W/>=7RW:NE4/8:aHL?,851[,YgG/CU:JY)8IcZEUPCT91UG7
:a9LXX>f:LT6?_H3(Y1K/F0.AMO0fS<6LA);]@+.5@I]&Ag[F/LDC&=P?L)e]QH_
PAFW38=JYHBCPLY2H>GFYb]5GIJIBI14<YgCD^0\f&S^-EW>RJ;<G[:e?N=@LXGU
EcQ_)XN[>T,L##>g<Le+O2D5fHJZG7Y=ZMZOYCV6(CD7b/IObZ;X@g+cd&-Ha_0d
ca2U^^VCE3ZeCFZKDX@QC@/I_f-Gc1Q<A<72OU;J:IO/d6:##;N9HEURd;,DLK4&
@bg=N^&1baa1<CPdRZbU,:fF7102W)P^4Y>_-LBT,OXYTN2>#EEPFa,eSF60LXZM
2(A[)P&L2[]9@)^2]U[1cf=&US+Gd.UE9Z:@(BS2ZM:.,J6_M+X-@9K?LA_C=@A_
RNQK5f24@3/gLbO-/G/Y38d1715PaPP#Bf@@eV5L,[7EGMAa:.K(]IdX)YQ:Zg3A
FL]_2[(.)WS864^SbefV6/e[):#:QEJ1cDL[S_Z8^WZNY6AbD@>((JRW#@Of\(A)
4ed5C^[SJ5.;WeQ+gMbN9I#33KSe0ZG,cNES?CL0LQdQY3KEKW9VdA&0OK9+[gN&
KF[M#BCf>A-&eHC@YSQS:9V#;6K3#:4(>L<A>47M>]KLW24@]71;XadcN.&67aXF
R7(M>C;[OE\4O];D3_aN<A/#MB.Eb=U6@((I4BGH:W[8EV^P9M8^+IO2;fOZM0V2
<T>:-@F^_\R^+_D9QDGTbGSO^B3EAYHFUJZg]-eUS;/E6_@7T+/Me&Q6=+^8[SP#
4caST([N;3.;Q_]8XW9F^:8bWNRcNAObMGbgPX&H&,P85^KNNW_@9c^^6ZZO1&J3
b<<e4g74:.Zg<R=]\K/Rf\DR30SUg/10Wcg8aC#BG&G<>cZF\6#fZGH4H,=&;P8U
XE@@FTDHC4R]DWJ[^T4J6B(IRO]V1(?NHTY6QC,-L3caK;e=VZEYDQ4.2EZXXCM-
HOd8fgg+,V6MPBAFU<#H9:(<^+)#OM1_L85G2.b,-Fd)4PIYeRPL=MK88;MT64eT
F:V-TKWdZ]SC<8.[Abdb/HVGQ7B(#QSf,R7bW]F5?1U21TLIQ#G[[&4PYG#d/a8D
Hc+d0DP4E<).@+JGV04bKIC-JL<ZQN@].bZ:3U@M@]72.f:aed_4E(V\UGfD4X&d
QKH:?0Nbd\&HY0XK+I-<N3/_ONXF21E?91P79G+V[3c^?;]YS8TgG[G#X^.e;&)d
a#4g04F96P9<JRaYNbRTS]0KF<A_EfB_ML0c^[D98?aFDbY=C0e^;OTNW+QGK3d+
@bA>HN;<ZUY^J,=ecW,HXWKP<[PRfM<^U@LFB>.V\V)bJ39.^_3GRF5e0^GDP5SO
eX5GJ>fN6HUTg,Ud1A2YI0V]-4bIc(??YUaM4(VC#J)gN0AI772YI3b@SJ=).O.:
Y4;050XFJZ<I4OY4D-SbOM5ESXVY5D<6Oef#RDL9bd?2N/Y(DOcG=[<EP.Y4d9?b
CD#N&cd]8RDCeNC-Yf061YV65J0JF0Q0)^X3C_K-)bGa#F5D?cWaC1_>18]WMaP=
Y)Ode.&<74-JK3?)7@8#D8-,RC1/N5ERN[6eW^1147KEgX/eFT-YH4d0V_WY[X2H
UX.@YA^?(S<MYL]A\g^HE;^Q9&DKe[&Q4MD\(K1f?=;S/JZ6BS6FBOKZK;(FD9DZ
_1F+3RRM-U@6]>NK;KA/3W@2fRR[AOG4]9VKK2+K[g:b1<)1Z0a9#bBW99g0f-NW
4feA23F/Z<>;^HK]1H_^#KT@9RS6[IJYH[fT/:3(<?/:NQHC-I/fCFK\;NDEJUaE
<a-O9^^/HWOf-(>2SUR/7N&RQ1;GLN6b#PTXZR,[FMJE7X69780EG]19.(T[6J.;
<.0QR(Q3.1(T-<=V:eSQU0VO9@-Ub1DNaLIC1?L=1#CFgKWFE<S=3RbY=UB1\MSE
<Q;L8JGC2.L42YEF_7Z2..O+A+Z8WCJW>20#dZFU9OKY0GXPO/K<>9f42ag:aD<;
544U4TM7O9S7AFHaC>c8)#1gTe1XI_V8Z3L#_9#;1_/?=YbG[XaG.N/;^&+@2BEN
K@7-ENA^TLE?[2(SD@_6,7dbIL2&RDJZX\-;URY6G]-G0OU\C37]P)_&3+Z]a1;7
e8]dPU+[[?&[L9)\>@a^ZE631.:K,Y.#SW9aKggb99:Z[-e_RBC\S5#Lf<2[F>d8
?Z-(;@.>ZIJ>X=/6)/Mb=#B-0?L?,:DXV@_>0e\S&L^A5(G>RX39#.WU2XN@/&0>
g2--.3Y[I0;#ba[;0#^fU\QC(B@CP=ZRC=B@;B5OgHN8SOeJ)DgZ9;f_[1@WHSA\
FHV14N_J_RCA8C^)IM1X])JfIQ4_?Hd/1<,<1NECEcf,f1>B1>9b.8\5P,((G\F3
N5]=ed@GDXdKY^DP.X0[@KTSFNT(Y@D.[.S+c5L2:U/O4eL)M#+=aNg^VJA:GN(#
d2S4GR94F\4=_+5?\&T2BXBd0+#_6T.?0J<a#aAQIf,NK][K&&5CT?@^-cHFSIDZ
JDKb7cGd1dB.UE[Bc4[Gb18Z1=eX1HB9SZe]\RdL-P&KNOIUYZKLg6EaGbgXU#<F
X9_2@Kd2JH/YD_=eK5/d,f1CFU44PNP7@4OB1DA8=S8g13IT9OQg:XJXf:#S0F9c
.:3]3JU8YKNc+dE(:NUDG:((^Kd2Z=F#RS)[[H1d9c?0[RTPZ^WaQDB0P^fTP>FQ
TG-a\UR,ZTI25++YEe:>.L+D:9eL#[5@(W^;\?^d_<.,>G6f6UGEQBOPJ)I;>b;)
AH=;FcX:\#?RfJ+B;10B;QO6OTQ-B(6KLY<5]7+5R/_=bfH7XJ@1K^=a:D)&V_X+
H&)WDeQ4+V6S281^5[L76=D04>:.fR0D+N@CG9+2]RE@8<e#/CbSNHWc>1)fIYP?
@7=6&PPQ1&KJ1UG91>aUNY50)df^.BN?#S-)^.7L9GJD@S[M3[6P>8O4c3YFX4BI
_gHc1]LOc57K=1g,24KdS>P4H/+#09B]&\-PXcQ2bgA^dFXD+aW3fLQe6SP/EK2Z
G/ca#P65OW)^:PTFZI>D8T6^7IHI3U.GESD^/Y(3?&5-J)26MPJ@H@0eU(;)L0Ra
CVAa_H]9)^2e7<.gLC7^GUc8a2W0NF.Y1-U\:L>]X1+\ZL06:e_e3Md^f]g:]\LE
NDJ+24fA>;9CE\=-d9R=g.@,KZ>5BX-c]DKBGbId@d5XCe6Z7=.3C9(HG9CK^2_f
7#D6</-BXHG[?0V?bB?,MTZ(I(OAV>S#Kg[TD.+T:ee?V=HVc/W8/]J7]AN_]f_F
f-\>;7I2)08EU)G=9)9,+,dL#Yc/P,YR6)?NLSSP92=&ADU3W8PSQPDF6R6N/QD;
@<7/_Tc1(^FR3^bZ)eF-;g@b=C;QD?]JBf0>DKV]Z9YGfC+P)Y.6fXeC<bCgU-XU
8#/C)I(8&GA&]>CJJWb-,fC(Z[PYS6QJd:_d^SURYFFUJAM9[Z.>:TdH[1]5bH^W
9Jc(9;e]Z.B+&Sd+/3AJ:.a31<,89RB5ML;R8,)SHGd0OWG@d3L/?:Pbd#A-IFMP
0BMFO\_[<cEBPEF?BKL&V)N0ZP(BR)OaE;EFLYg5KSeY8144\#J[C/@X?eb6.R+D
Y984gX2P=U9KYOY75W6M[BaWdTM4MXC2PWK-?^8.7<++9cF8LN:6=LYL/LF<=[BG
5Gf;9?]C?U1S8eadUP=4;=Ha>EK&4#+]Y2UMWC;SFE,+Q?F^#.fWH5aKFJ42\R2;
1[C//,=\0<027VI+(/]/<I#=gR<_U:.9@RO]b=/OK[88a(7EaF.HR<6+1fVME]B.
\dEfGPE??8@EW=4&Z-,(?V+#+0E0^1:9),[QU\253).O#5A]AN5)3@7g+/DH.&&^
1_QE?TP<XP:fN[6:U1@S^^aA?c/;W);W9CO1F-7@#Ra\4N688&[3V3D@P#J2-58?
&H>^8B]\HUH+SYU9\[[^cEGaHRc;:^2VFANF1TY9>#WPc\fNY[PeI.-/:Ya7Pa^C
?SDIcB1LD==6:&PVK]J\#EW(3+]4Q+:dCK8Ob@/KdB<BD@Vc58LFPVY1929V=O#R
bP<gU2^4\;)g22dL1d>(eQXbA?W)@T?1KH3WWKTQ1e1-QeJ/gNVS4,QE8O:FWI[#
Kg),g(O^KH#,>]c.6#FH+\=IDf8N-#\#F/>4T>2(3BNE>/T#S?8bVWHWU1S<64^]
<)Z4&W>M@9)8NCZ=b3G]O[8HJf_0E,9.<K/\:3(#[g=H#RG?S//>aX5.IQS+e^5V
B^(e4eFbLGIP?da+O@0Ja^=L/b>9eF&bcd78:QaeIZH/>HBXN]fUT.2JWDOCW/_W
<be:2&.^^=(N8.8E3W5_^CQTg_fN@7+ZR/3I7Hb63E;2.Z0fMXOXP^D=R-84RUUW
2JKNCPZbJLfE?K@0T?-2^\@7<QI\POH8ED22ISWQ5IHY@Q@K_EY;HK2I#WX0V1d=
0\1JXO?O.GYMS2e\fG(_EVgVY2<&ZL,EM[=AW\](0(YW#GF1b21VOYH]5+aL#Ob0
5(EZJM?-2@L^]TN>dA,(bC3U^D0d+6HV6A[\cB1CT,\[T)M3U@,0GJJD64Fd/dQ7
M5WY&UG,?d:1ca&[C#LBR\.OL9)2H(VYAGZDLdOS:XD^dOYAH44EH_aF59>8H#G+
2=7-dFaCQ/dP80DP(+a.eXNc4W4DJXS_;eU?Y3_W:].ERVN]RZC94R?\A<aX?Ne5
._:[CV9=WcU[K)M2fY??_\b-)d;ODW0efe9KBAK5LSLAEN>W)N@E(4(dMQ3D6d33
HcD2\(9<+bVBR,UF->.^bL..TBI6]T4Sg(H=<Vb.;NQV5F5N@RaB2]BX9OM)34(.
;FL9fR[(6#NFZ9,fY3]FaS[=]&Of:[QA;:TA4YcJURPIa(Qa9^gZ7c=V6RK7C-PE
C;@2R-eg=JBMJC^G.bZ\EW,cU=K;b@e\9F]RSDC^=V\Ngg:30K0NN;C:fI(b/XNA
[?.,@,(GVUX.R.R[0D^=WRDRQ&K2^3dSe#\I>Lc;:J6MTL(M&0>UD9^KR8<\cHO^
42JQOKHgD_PBYd?TN5[MQP/S5U0M,X)<(#P=_1+A+Q9U^;aA;,DfQCAA3+O;IRVT
H,Td#>O@QYR?d<J/_9E#D7VT3/8,&TS6:U4;3V&B,K1]S_6G,Ve=\2H^ULc,^U.9
_NJF;a?,6ST[M2.b7WI/67(\cgGEgO@D[T-)f1?<#e@DJNJ4UBDJ@bY;_ZBS@(2J
/#UCN&&S/\-E+XD4@4D_\eW]3M>LdeG@><VYbS,DcgF7.<[gF>6G4YVOP:>O=\V0
T)ALVXgReGZ^-PbgW/P4T^49Rb.1C><>K3W.C2M)>)RQ=bHXaI:bM-UQP5PB0/fH
M\[_4g\E<d4?GcCVN6AcSeQ3UOEQL5)7[CCC]4_GCaBP.f75@FKdCB<V2_C.77Qe
H#XRb:Q8^+8H##:V/D1@Q,Z_+7S6Y>f[b:HA\3@(fD#&Ib#DT.^@\PXQeb.6[4/M
caVS:=EEW?E5H_8KF7,V]A=M+gZb/U-b/_F<5G^CfAM-GZ>FDV6[[K=-_(]AfGJ/
D4CT447X-&1?8R_X/\1c5N@36@(.Y1FEN6f=_;f/.=MHRO/<ED_;UH9H\6]X3:@.
a2YZZc<(6/>58-WNAf\WCOK\KXa9/,Ze+KM5HKV,X>[FDC/]N_\2/X38&VDD/5Va
^;()0G0Hcc)<D0VERO#4?O#<=Wf0X31b@-=XOb,We.-\d=5c_Ae4Rg=<=GeYa^:A
FHQ(e#GCHP(&C#Qg1cZW?;3^H+TGa?<H)RTIG,3/CV]c)MKgB/CTUPI0M_]=6:JH
CTPU=(\ZP.3Va0XZ_3dF\WQ4aXYaEaMU;D6f#LRgQ0_EWJ@Yf33f5gFKN2D1gH&J
E/LQO<^@C>&;cZCd&0Cc,MQ_B5?U/(EA25#J2\W_(I05c4TR3bI_-#df&XG&.g:M
S9MJ:D,LM1>4J63DW+,PV60I?2<T1;DZTBVE(I\3+OS9:?&MM#JaFWSX@C9?_GXH
7=SPS.H^\Od>_d4<&O&7=([2e5:AAfTHO.?IKY/N5:KA33bI17XR;7c.9M.F1=YJ
2;KK6gefKe>VN:cc[G;Sd?665])QIK6g7:_A_LJR84Kfe2,,JERJP1:86UVD_(LS
#1UgU)0E2Kf#Aca=AE&M<C^g]F]6&C=XY8Y80_Yb#0#Ag7-@K:WTE?aSaB2ZcO<g
@eMcNN-<,Gc?(F4_B/>MA(?-,(.3IRDP]KIf/?B#W.ZK1:\a(C+@X<e1g9Z@a3V4
C[>CBPO#.NOAJ.[&X1#UI^_Kbc-6<19Y+1U;B]Jb/1]/aJ#LeMB./239d#(X\gC)
8LaIRdHJC.K+ZWC3dE3/D4TTJdDX(@,ME1_/+MD7I,VANG?JceNd93#+.,G+Fe:#
g/0NKPXW)Ve[f#R:Bd#WNIc3/IWM]>4A556<C=+3AOd(aCJ0@bHg#:84C2gb@E:M
7K[2J9^(dI4c1UM7.AH^T[P,/VF,+g<J\aY\fWYPT50]b1+LJe4YQZ#F@GRB+/e_
+_E6:Q>dPeb)0NUL\698edBG]C2^P,bFLdUL.2^/;?eIUNK_AbO8c])c6.E6N1T3
;FDU)1e5.b-V:Fa+.IS1;_dX;V.)<HD8TGUPW=36R-0&<OTT4M7g#a[E0AR)XU@@
+XgYH=UYTJ&f-fEMLB2B+M>=Ic(fQKV@2=8^O>^H==.9<0Qd@4X)C.,Q:Z]EXVgN
=&MKL&G]@+\#V6-.?B;aQE#NK569\A]SH@1A8+Z(P2(Q>9^RDNS3egeB3\->5BW9
7P5g2U,PX&@9)H>(E-U_^2G9_:bZE9_e\4gG/52K\JNL9X7Oc)P>1::,YF.8,8gH
#WP=#a?[.8HS293Z]_^)2J,)ZFJ;A4]c/R#L:Y]^C.eAO>ZX4:R7@S[N+fFD-:44
TbQLK7)FVJS@Y6W[1\XKa>-)&G_\b<+c@L3FKNZBK3.G\Cf9UT9E6+Q(+=NI?5,6
4.PVZ:LJ-?)]J[[;1Xc&N5E1-Y+O5I))))-,>/G#3LV1CGNN7GKL0F;^;]^g.#14
0+Xe1#/1QL2>I<&K(Df[O_/7f>fF)aSZ0b<W\H7b=IYHP#9D9(;[4?IV6C7e&:=D
M(g^;V@L#G.5.0]JCY<gOR1ZKXA^;/[WXf979W;eK\8YA=.8/eN[8NfB3gQZQ.\Z
0gJ3JWUcdX5P(^Xc9_DU22C\F9]Ib1=PbI;HSLG)WW#6f?6Ef]/\\]fY,IR@K1]Q
Q9_L#V\CG(F#fL2/1DUAKY&]fERH_0FCG_V\(9bSKdGb>[Y>3TI7X24;8OB);b18
b^ZC1Mg8[/C6A_VZaXBe_^Qd194@G:fb\SM]<.FZL?E\S;#,11dUKbE/[+BI#06O
3<U]+XKDAS:36L>]eV,fSI7BNf/gYKWWE[YV&c[;81>(F(c\X7U_)53:ZV-,769C
4:dJ^\Y(HQ/^JXP\5@I2AS++eTG-7>J@FC2D(PKJdS4bC:)K0O:VLOD__^UB70D>
Y;CFJa_/TGLNW/S&A3P+[:b6&61e_Ne0=24Y-))0&9E\(@#6#cOJ59dQ1V\Q<9)V
0b2DD.5NB>P5L5C/3Wfg[c.#+d-2RE=RecJeJ^@UcM&ZQ\Gbe)M^46<)NWDTJ8E]
.8MB/H)4RYgW8/Y?Be^CW1BOa[283Je-27:KB[/6A(+X\MDU[HO^FgbZc)4TO.2;
X]-c/J,PJc7+^_CSVcN^5Z+KLSdZS>8:B/gIQ>W0,KS8/S5C56SS5OAJLfb3<Y3>
[4.@\gCa<I[.BQ/1e)?T&4cLdg,b\-9eGW/-Y2P;>)Ge<XI-@Q#V^9fY9e4YBG[B
(:H3FL85\:]/AQ@eeF,Yc8V,+@^W0a)=F]+HNc2@7cAN\cOW1e9_Gd^XW/IH9.cQ
MG35_a@f[>64dT3YWI&?O7<?@cDaQ;OF2c.OOc9M6_;Vd0GT2]5I([dS\0N=W0d(
R^:1@cN-(.UV=OA[,A:EC6>>0:66^#:c3:=(HSY0TQAeC+97__aGJD&&M<63UDb3
T4,Mg/U;8bc.06ZY0[3U+FHE5Y01DJ^W<Md2+Q2&:I87SF;FZcOBM]I[+6<-cKZO
8:@e?^)+],9I?)DRF1.VT@>M]@2Vf,=RdKJ(=EA]ET0LQLFNSPER1AV^_M5>A1,N
:6NIAIP3B&AOU.d=Bbd\\\+A4TJW\4;XO/]#5)H3/@^1PKdR1TD-g-)aN1Wf&.2I
#)[I:][ELgf.d#N:W__bWe@#]^((1;R+27&>;73KUR(D/f@:Y&I96.b0Q_V<#gX)
4R(E6)9V)4#XG048#G4eH<XNF>_TQD29VR;)4d0R0?O,AV2UEZ>/(-b_3-MUeYIL
#d@:e:Q3a4OLHfL=KZ<=&FYae7-ZL.0XRM8fd;Z5We\457\PVg>Y^)cd/fdceSUb
5d=BLDBd9:XE@5RY^_9#)-2,OGTJ?6V7&[T,2c35DBf[f(80YCRT<Mf0Lb[\e&VU
WY_NdR0K58\=<@Pa@Ag-2-?_e(1.F0G7,0(?d>+Z+I7+;26Ubf2][#Z^L@9JMTVa
1W<E[]FT\SUN2@]ORLeW;3F2?.CE<D>5Z]KO4?TVP2bN-KXP[fg.e@#[;-N:7V?<
Y9M-C??7IOPEWP1)3VS1<)GO:<ECM#7#8WEDW8\R6UaL28][W<2F,EV>&05XV=::
0FR+-FJIG1RSK_^O>2V@:5A2Ld<3a[,^KBScC#NN2;,=]?5B9BWZ@MW6+6bH6[];
eX5U7^7Aa6NSYbLAbQUa<N2La6F^Qf\XeZGRcJcX;;UZLZ\;W7dB,0FaeSCTR=_c
b?-H:,V#V<,L=TA8<&-EdbSBdTNJOHB7c7D[a+E9+4C02QYSYOCW[HaMDH5_X-LO
:V42cOcPCaI/[YPdN)HEV.N-e.DN-RK[B7cW2aaU.#MSFRWH-_P7dCHe6V=8BS[6
UE6PSQJ=895BS_&>+])K1SIB)J:&gNC+;()#R-A^e@EA)7bc].f84W3B=[7b07L;
0Q]=J:dVS4<<5BX9=FR.aE8C90:DO)2R5)B9:[:Sa>a)POSWaZVBDD(;8Z8GL[^[
Z5^D_g.&KJJ9&GR\(-4Y-@ZcQ.(ROJ3ZBf#[-+T_d1RP:<64cD/ZWL[,)KE,c3<b
HRE>OZ](e^/VS\/5/a7-\V]A4ZDcIgTI9E)7.B<1IQ6?+DSEN-USSS/P?.e2=:Ld
T7&81S0eM1^]>#^#,++S.]I2@0JB)YBO.f9V=5&C\_M1(S,&2.]?0-1@OH>TM<f4
5E/#fBM;HXQFA+c9<^,UI_2)Y<XWbL6D/FDZL-0J/RU+6<75-&VRBV]=aWH0^Z;2
YVD[>c>\S<10DK9VdE2I,VaM#0>816+7T#-[g>.HP9)+f#()]2\]MR][RdS,(NBH
EP8[KE8ES3-N;-2V@fdQB<IEaC[2c#.WQeAfDNDNWQL=>[&ZE/:+?/C6bQ;2Q+D&
NbH/X,?/-Y,;1a;cN#BB#,e08>JK;+cOOU/V2YJg5d4)1Y)JONIG&Of.2YVUbJ51
SV^\(R9Z:T:[g0,SER56Wa?U=[K?Y8)Bca3RgVU#H+(c.&KR65QC6<5_SP/_0]&/
;XNaN.MFIfARN;)A)7e9#Lg]7g0Z1Lf0GIZd_FbeV+Q[)<KM_cJHD9g@X-,F86;;
=#83D^O^VAOOV-+G:+H3-GI0Rc.fXGaK._-&<gH60U5.YOO5Q@5?#eGDW];f;fa/
60BT&J?C3IO_L/394>dKXZG@[_fG87TS^,S5.9L8@f5X3##_>MV6A/-6_YZW9=Rb
?8#T@J\W:aEQM[e1).g-;CbAXH7#KNL;]g(<faSE<JFff[VLXWW\^,A6f88E+7Cg
0cNMe8Xd(eQdL69GDQ.Dd?1/_3a7+LH:1N3fMZ+[,^JMEE^56T#_U9UUgP@J6[09
fT)^WA;a0fU(Df1HZfedB@X754R,EaZV>]Ub.@JMSZSTIGX4D4f/U_E(E6XV7;1Z
T#Z.bYY:\7BB?ZNTN>M\+MZGgM?egV0FS?d<0MLT:f.CO[UERPOgD8gQ@JBY0O9.
1@P-.99;>&E0fK>:&#:FT(<<@K6DU1JRRO3EC-SJ;7:I1#@D1d8U(YB:@\=Jd((0
/1LD12gI)7US=GPSBC7bNIZ#S+T-Q\<G;]EPBZ?Q?2[4T2Z=Y(TZ9V\LUPY8?AD3
ULHgOORE0BeSZ;9?>Y^2KZ4[=,O];BQM-9C<+3-Pf#I]S0B28[5_I/4\Q6_@CIQ>
H^LcU5K>MU5MR(Qe__>:(>5^4@BVf=A1&,,C0INcX\XWR,O(T9;MMIL<1P^Ae-C=
.1DVO]EIWO_eA4RC#Q4,^^=bFP]&<196;\A(JGY^QD#,45)]^<\3I10,Db4+-C3<
>CfFT:@N=-W#LA+6HZZR=PM#;,=NA+;I+bU;C_4SJ121O[4J:5Q6M]W.6KZ(8+@2
D3HM63<=_+GMT0L-QDKR.8cWJ@JDc5EAV_M20OM?JH]N,]WNgH54dZcGG^,OG3^]
;#8<BB2:gG+@N7\.=6VcLM-9@;,)\H9.11C/,@JUcF,&9\199VLK6(U^ab^;>;HO
fM(g3gQUN+L^T96ARd^(H48^6P9](]OJ1S6W_2Y,:@9ea1\N]0Y05+/=B&N=:gd:
:TQ&B3Yb;;aVPbPW]gP,89^3:M&:B4-RcPfg@I/_G]CQ)DVZ\)+D(6(AE,g64C5V
5Ca5.4:R=&8gA/O^S1P[M@O@Mc1N:[g^,>O35LD74=8c</9UN_@HQ7TQ2cLP@]<F
W5R05eLX(=dGR,^0+_\LHGN:TeCgfQLWXgL)P)EHEOSL/1-Z5_8.)F1/]b1KY?bb
8+-H=_J#_5:(LO1Q\U/4Nc^e]&/Y^e>=g6JZ[I7cRA+MfcA^,E/[0-AD^8(X9+eb
OJ7U#B@5\JOP;0bM9]2A/J<Yg,P-d:38KccOT\P82LBYSOeZA6IGI1.fBTceSFB)
V)DXXa:^)/)PKffZdH+:M.(&J/]M9PA[K#Eb?WL^752N8C9/W9ZN^8R)Kbc].+aL
/33_;0TY=WA+@#FFc\b@X9RJFM\c/SNZE-?8PaZZeeIaDb\cKVDaZ4R80F0:^^?N
bU[?QeSGG_A/Jg8-cJ#V059JQKPEaa)f6D<e.A51.Z8a<P#R43>)7)D;LQU8E02X
P>L\(JVF6d?02;ICY5(S\LVd7,AL_PBX4b^K4-.d/W@/JSRg<.86SMf#QFUc^5]4
FHgT9PP:QSCD.Pc2-WRHZOgP]UDKGf:WFDXZ9&I2#^^4@FV<EU6T_@)88NT>f=:&
Z:2H=\bQ]3D=OX8ceV;\0O_TgbFDJOX3+P-[>01MNg2^,J8?eJaI>cN>ZJ-TT])<
&6Xf89Re8DSVgO\GPRZ@I6PPSFA@::8-?Jdg,R^IG52X5V^[1U90NFH3/+;#e6H#
C8>f[]SHfK9LFMd6aYTU+P\<B4fGd0J3J>67E7?N27=&@?NS>B.@XSeSgGRY]TId
F1:[2Bgb^]Fd7F&AC2-(ec>RH1-bfT-\J&?2PN]YR;?7(&BZA6.:aV(gfP0[[7F7
/UIZEb1H8I0;R7g8GYIR4ggggP@.A@f_A3JJ<,)43NZUP7\:eUU))6?:TZ;BZ7EO
A(7#BKYKBGX-Yd_H0TAE4/\YTeRef,-bMF#CXBF;<0F/GMcB+HG?3^d>#D)4>#M6
?a-/B/TBO.,-ac5B08]D37gCY6UTGT;f:8BA0U:D@HF_X9IKL^Uaf8,KN:A?,UMG
C7X[Z\I,>UJ6CPMg)O1;(A&1[,PZKPICK1dSa2.\FKU_.T9;\H]N(<4\0H9/7Q&M
WA;CIOKMIa5\<A+TJIFGS8Q\#cP@X4)[(KEF\KR>)&V1,&Pd,@34W.[<0^8=RNdJ
BGG>EYX+cOO^K#U_HaZBXPB/#HZR.+T7dT;[EWHA;Rc35)58PB).GPJc;-O-_g85
d@YIUOaSA^<4PAd@c&NANX>T;O+a#.RY15F95)^a&[d)8NGbYaaDf.WDfV?2aG02
ICa/(T\+7:OGP,EGM,EDW:#C+CP>BH9NH]QGDD66>?)JC?559(3SMT[MTX\7ZGFU
<BLQe]=0Za(L\F@ZRMAb/YI2Z@4RE#Y>N./DVC)VRJP(S>U3CE.b:D5.3IX._=&\
eC&Gc:J,>d;0,<?Nb[._-?3>VXdI>TX5B5H#EYOA]b?\g4:KZZ]f&e#_X>9;F0&\
0M@&9TQ5gB7IJf:7d;@=?+/8OV#LUL\M>c8(PW2PPVKTcZ8V-E=(<^,RCA)H@NU.
G>gJC^_JYVEL,Z0/];D^<F#9),WUGHWD[S;Z^XKEFCD()eAfWH-K>7QW(-;BH\97
=T/V9/2H26S-S[E=.6NPg5Gge/I\/B>S3Q8e.=F1F(OFAG_F)C8cPY:fIO(LMG.S
>JeMZC<R2;0d47>\]-OAKcaKTLR+c;B+CI[);O42g#]4DeUMHKR_;1OWO3[d(Z??
^dU^3)c21R0.U]]GgR^\3N85PaCaHfMCU507QCP>Z\OF,eM44SfK5B86.bL1LGKY
eGf2CaRL\Z<cMML@W<Q1.]9ASb&\^.);U4Z>;cbU6Y52S<]6+?#=LOa8H@g2(9d^
+II5^K>3J??/E;2;_\0b;;_gC;/R[#L;_c)S>b,383Z07Y_K4Z,JT7Z?,,-SeBW2
WagOQ?d<Ab[db(X+1c)&TTU(>3(^Sc2H27SE&F4<AbEe#\X1E5ZK>1NeY&fT7H-<
aO_7H_.@N;91E?PJ8AK50QY).3NW.#42?63-6N/XWN#NM][#J5V.UD@87^eAfe5)
L[#Y#3Xd6X=N?ebL5Q?Oc8M@SCbbP\X#^)7ZaN;SK>;B9bCa9W,Wg.^?-(,c]DLG
4:C[K0@EZBOe+.7Q-3B,DT-C?SB8f)KS\M-[[/7fN_2E9MJHOC=b?G-S;:_+SAM8
NFI[fU0:0a&?fQT6R=5X5H8L265(H,;V]3NU^e.>SEE_X7#VbNW-c&:)OKQWI9S(
.a>_H(I2gUEVZ0S4^U7Qb8:)CPTAA]RR[6R.g=UONY8OCA_1V;?M6WGWEPa?#]\.
:0Z#_T[)fed(/4._D27W-JQAPT&8AeA^;<Y94eO<L^Z5=cE:)YXI8\35MVaIfVHR
cSbS<([F24P6.]Le#gL-MH8Dga.;^J8.fKV6H_3\0d?>SA.B4b7@=<.A95E_PW_8
<DQ.R^L5X^OBRB]=)KD\H&H6YON717\Z^&WBK.OQKc.f\90f;/67ML]J<:MFI+^f
RKc:SNAJb1)YC80bbW(R0cc0J03/cf)\AefPFG/MIXV6)[be3dNPbA)aT(B\7T2c
fXV7a.+g;_f&TIT(IB:ZDDG70;C@\c4>4Qe_#_P^\GPR\PQU4,g9>[C(G@2D_@84
>QZe2?@;[&NCFO&1WA[/Q\U:>4CW]##8)0.[78b^O&L4JG=QRBR+g(6aV24D]G,\
G#J5OPWBH1F1H)5/:e+5Q9]ER&14gEVS=@Kg\b_BC6)QC3=7M8XJFPP5abT@(1_Z
W=VW-\A)6^-H92XHZ]87L&P@E?UCPbD:LD-,XK#0J?&:EBL^A69PbaHE9&Z)WP(Y
85C6+1@E[a(_=QX:4VUQ16TPKRK8FE7@g^&3)Q(WB1JIAHTeJ;fW5V.TU3X5=&BM
OP\6&9HFbb3A5[ZW._4XM55W1E98D^>+MXWc;E.L4daP7+SaHd19=#?H6L?=e&W8
CB#.TEJ;O(X,QKI.P2R-PT<//IBC4@Y&d1GI2F71^FP,=g<PFGZ0MNU9Pg..<da[
0+>=>I8##N2\6eg^D0EegGC7JF9XgW:4a5fV)ca2V2:-3DaUINCe;):/YC<9Sb,A
WY08f>.L,YX]C(Q8.bW=]6<6K@OQL6I]BPGc4Z7;dcd7&>L=(>gV+<(ET.J7b/SM
RRR)]\eQSb<8S6[VcfcK7^#d5EGce4+b/=P/)G,5ST)4d&ADdb)TM23E^&.R3C3@
5g<MMNY^(C1LX434dF7#35@MSg8e,Rb^]R.4dG9HIG&3J?(4IQ=4)BIb53gQO(TS
==:0PHa,I?:.)+5KEI+cJKMH+_fKM@=)OLO:,g>4c;=d4Le6FZd6B,]_G(TC.EKF
e\6_WDRbGYeg>9,RLeO@N15<Q\8)\ETI1?dO@;5\>D6Q8[4QP__OSB3ZB-D-ag.+
@-_aMQ4_VZA1FdAU:PP.JS_NB./2NJC_>A3LTQ:0PNR<a6D3gI_O18?e2f?MebV<
>EY/W;=#gEJ,4[SQY@/V#U=e84KS3K>:^_^KfB2bM,KCf22/4CWe#B1BY=gQ#<M9
:F-AWDE/&4R1:5:^[M+:_X-;]8_0aB49O5USZ,LfJ4YWAKU=f&aC/LBQKD,fMO/W
Q34K<1bOBE^,GK&MA+-f7I?V=2>a0,d;IcF:,HW;KN+-U8g#6)C7FaLL:SdFNNDe
Y.EG=-[O=ZH-\XK.UR6#YA#-)FdTNC(JY5ZJ1FL<QEKB/KZ^2.ZIVD#M<aU(MaWJ
eVY9P>J3@WEa[BNXO3f&/H1,0T26P@/3>=Y@27N#<g]1F>A)&N(--PMg=FV+;,)f
WEP1A:GSZBXDRV_2T>IF2^?-6L&MU7YG8dRX[]Z2c#cHEGcL912eN4.OJP8\8[EL
H9(16LJRO9LEHaeVd7;M[KU]FU379W^UGXX>_4?SQ,)6;K4<6JGdU<)RC#7D?b=[
(bHW#dcJ^Ta26<N^#0Y;d8]3,VKL_+dRd79Z/&dJ?5cUCBWZaNV[UP8dP&2.&IEY
07<2E;UGVTTY1XDRTNAXNFWcHD/Y^(#,R[e2bP8bZ6c8)H\bgN4_VT3=^FZ7WeFS
8X8c/[^G3??SN6.NW8[;a&7dN#(T85PFfFPV1XQUPHYHBK<K+GX#>g/c&dYf]L+C
AJC58.&9cU3fYV<d?cW&df2_18&[f,=#A)T](/6TKQ<g:?-2b=;CRZeTR0AHI@XF
#L<aCGdMK39fCG,g/A<E>7PHfNf3R,GL.e;H@:]-Q_I0c<HRdWe-cU,HffN,_F38
,R9O5G.V+>U]CR9M<;baMC5Be&34WPWcZ1EcR3<X>fMT3SV^P5-+CV[3,K(ecaUe
g2b(V41JL[KD,:FSPNV_XT)3K(D\ZUX>YcYG?2(]5EPY-V]_FNaVX29M#Y.EE5^B
AP7d\aaK=4:NA;^@gCg#K[JBg)<?+Df7I_?V3LKD&[^bH=c.R=g52@TKQV#J>7\L
D6,&gL2)(]_3cdST(.&NO7CEG/B,^g[RGE]_DJ/V1D,Adf^PD-+g8FG-@/OISG<M
ZFaGO_GND2)FM+fRX:H=69Q+[3ddDPe;Rd/;/9J0F6Y2dUP-[0BP9U:E>=QUON\,
LO_[GH)SV5>P#,XPN;)\A===aQ>ZH2)af)4X^PeZ#H()+]19UF90;f7b?ABWW:KC
Y)WRA.BV/Y&Z,ZQ_#)AEWB<E>aLOR#[#WV\A4(A./B-7d)Y@afSKWN\0T:+gb\VI
29^HTDD<(XE(,@#ePg5a)EFb)/Gf=RH+UbcG&7NF5^Cf#](U7#+>DW5A.CIN040\
9.4LKOQNV,+1(U^M4b8G<>HGTSC]9.aC4XZ5gb).))WA)K9(NL]T@K-YaG/][?CL
)ODCSU,OH+2.57,8(@a86\//&V6X6C\CVMaUZ6TfOe^B+e8)ab(]?,D,ME(c=Q@^
G/F8^9dO4ME?ETaeQV1J]7^VTH[e\:Z^(\<U9LdcK)3KdG(7(?Z1TgK7HZa><7P.
QUYXHIS]Y1f#U2J/f#J<8D4>[bae-BYM;V/NTOJNLGN6AfZT(\N]@Rg(Y-Zb:ML&
K:H/?dY#Z;EBE]YcLK>DHR+2K/7TE2]M]Bb=]4-+>ZNHb.ROSKU8:[JS(e/+BGME
@/LQVP#->(\DT#AD2c]e30#;[ZENa8^/VX,FL_)f1a.eZM42(@fFI>#/GfWL?:[3
.MF^0gE^3>\S=XOE--9dWg2P]5X9E..B:E.\_g<03GaOTfHNDKO\FF9-T>Q1D;--
8IPT37c>/S4g\D;aa3GC2U@]GM(eCf&)>&G7GDBM&B0AWPCMXP-B.Wf^A-QcQW(Q
)Ob5RGNP4d.U5U<[I4I;Tf6BDX1g4f,(KDb5]^L.#4-=XDSK0B.<aX-EA3DLRW9H
MQ]DO8THScV>K9F8S#DS=aWNG=]\-.0CbM.0A=K6?/E.agSfX)2PH;K3E73D);CT
[2LTc/cYUZ_/d?CdSGTa0G/W.M3[<-,/@4TAQ.cda+1QfA,@J:cd4aO\Gc&&ga:O
:AU2BNe,-S)K9O,+e&dH<=CIJ49fGH#/BZ-bYfAYW@9-X81#_[KM6^eV/>g]9JMZ
#?If5C&?@ZJQ\-+23WbgOHJfAOENe&QgZU:5/?5]@#fPY;TO-(@;E:<@L>Wcb9+[
EB51O)e\Ba,^<A6,.,\LW8<AZOH/@e\&_DCR<TU^eOOU#W(74g(e6#f>3<QYg_Y4
#JXJO(b?V+HUQE5L=JZX2gS;,<NPT[RMc_b3NEEQHb@CE]A&3e0f12RTJePdLa5b
9V6f/-bO&9bAfYK]2_)e+7&4_Y[>N?4V3KC2-HW01=Wd)a0)ZSN17B.a]I_.9+<G
I&SZ^JG5S:-CUUHaFY\g/.7;U:M3.C#M\#RQFeT84]RgPOU-+0\:;YO6+4JLCM1B
4809>PN_<VZeL^Y6=VBW0+B^^I^04M8JY/TF06I1+X<HLgN#KG]W<2/_59\V@SQ?
JgCFe3cWK6cIIfY]d/6WHXE(a.=M/MM@^C3OQ\d:5H(DZ7,#>3TQ\)5&8(L8F63_
K.FAGX1UZ;M2EW;/E/W.H2E(5$
`endprotected
endmodule