//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2025 ICLAB FALL Course
//   Lab08       : Testbench and Pattern
//   Author      : Ying-Yu (Inyi) Wang
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : v4.0
//   Note : PATTERN w/o CG
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################



module PATTERN
`protected
7..<@GXN9YF>/M?d97D:13Q^d,gC5:^(6+8,ACMPcU++bC9[>?Z8+)..G]<Jd.G4
a4Y#c<a,L>O[\WTgMN60eXg98Z<g23Zc7#)P7=F(AJ8JB^-YEg+:OOM4,-4X1\8Z
0?A3NSRC&>b.IPebV+98cH;#DGKJcR&8Ua2AEP[U,&KDDUe&74DM,5(ZQES,YEG=
6cb&,I\._P8C>LK)H.:4YDB/.NQR>IS0?:JLM^)^=H/(-/A/<4/ARV<FW_@TX(MY
(MSKbT@^ZfRJd<S?<E&N7QD5=B/5XPS>22F5]ZE(+NUF/#\#a2]@eGI;eZ\c>\>L
A>J(9T_;CGfMaYYT+[]=[Ta@4ZOT]H(WN>I<dLYa48J;^YC1b9J;XB@;ISbPe]AU
]bC3-_Yc;DPP.4NgW^D&J]L2\R?3T(81-f@#AJN_Fa3dY?NI/K(],,(;7]&T3ZI]
CdR\HK-(+=CT>b=b^JARg7@TE)=OSZPCbf9Xd@STe\FT06Q0IB-E0D>?^e;9e@F8
<28c3#COcAPSc7C)N)ZJV0?KG55.aFbO;L3Abe7A&8/SK-V.a#.=M:D9IE9e5T],
d@V^fC(.8O_3A01Y(=6@;X_IU<>Pb[HGb?+(bTa@,SKg_A@A42f+XOb9;,M.d1K6
<L2UH:QMg?,FQH,=38LeIP>c<0Q#eV-T_G^Q9f(Sd0-_A,AA-^>>fGDQGY(<>D..
2W=F5T^/,@)g_AS^(BAc4NO#VTB4dP=/S#TQC;8#0Gf:e+Z<M>_6d>;KU)2aKER)
WX?NYPB2VXTDGUW@P-_[?KR@5FN9G78>6Q7-GU<P4)QVac(53=d=Mc33b4M63302
TGBR@[(6TO<:]f9Q4fb;d_8U@=fda<#YNcO]?UB[(?U=BJJ7E.5)-0;QNdJ[AH5R
4ZPA6XV5T8-<CB9.d^XDTPZ6?MfagK+b1F9XNb.]59&A6RC>_/?+0\PeY9Y42XRV
<c^U/0__C+e2C-H:W[7VYM:Z>_]I_<F@@ZcVN9M;R5++C#-eTaaT_[b,G6a]7_M=
VNNM?f&C2^GJ6YCT#6V:\R41:/5TEP:JBe]2F]+@D5BW+X?@Vf]HI(A1UL:KdZ/Z
Bc&=Xc9ZHM<c4Q8ZHK/5Mf3V>P97YZ>W,bOTV)T(J4Ce43O\/CU>N5S^=dH;]#)?
BBHKGQI(AF86HC7FRZ<XR_+0^FJ+6C.@-]1COD@e7f2:;9#2?Jc([eKA4EGL@IM8
T+F-;IE@Z(cR),_6[1B\I)]g0Z6R695YR-<(E=&Qc2PF0d9GW0+B5aE=+#[M+<(g
PQBLH=&6T/.1WF+JWX3P@V,gH9:++=10dRY-0WI-G7NJ@V3&J]S]>)QX60D-QK.b
MKXIS(B5/#QX9-?PWV\FSY[,Tc\#[3KEU=X_dCP1ATTERX#LJ?Q_SH>3A]V6[+f;
MU:&AQ97I9(>e:.<g=[6#/+Q@8GQ]2I?-+3<DM&DARY&[@@G_[Z?-=LG4gK2K>Af
8F-c&FA9F]]RP_^^L^Y[Q:d7S84UN5-_<8]cK/[RX?f5MK/cHC@6R5NH8fR&OXR7
2.5=\VC[)J_&FZ=#>FBKY&O20TBgF[/CYS=?+/L[]EWQ0GG#7UI+&W2d]O8\WVf&
,UEX>?X/Z_IK)\O.97Q^WB:-R77Y<S&8?42-;L@T7D9Wb(,3C@b2CGddJFAS<ZSb
)X_Ngcd(Qe_geLZeH^fPZ=^7BF,_><:^O10_1[/NA8EP,-OJHbHW3Se33X0H7:1M
Z^CZ:Zbb759Q2QTe].?Ag1:F[MVB6&;KTcD,I@2;fc)TZBR&2&Fb623RY=?0WG6D
<F#=?2G#bd.A3g2NL3b/f0[9LF:LdN]VGbPZ-g34HS30S@:7()BReO4cGH9_(76(
WXUVeG/FbC6:#J\V@2Y0BNPGa.Ua6c.Cd1XI/&@6>763V.[^G:E8,K@KFW6J8N[.
@:d5]NN\d+\2NY8LYKIYQg@=C2IJYe]99S[?[8Z:_aLd[a[26MWC)Ge2UF=d<:?5
MgYN//V8+2cYK#(SD_&g>W.^4BJX7I))Da>NX=A)-fT/bQf3,CW/N:DZbUD3)\PX
EEJg_eN-<@>gT?SXQgGL722dMQ[<\8IY7PLF>S6eXH>VJ]M&E7/L]-GDQTEd3MK)
WU2/FHc&JH=2U>Tf7gdK9;C,IgP;G1cM/SHYBF&.Q^R_aY?@#?^8=bCR3K0G;2@F
D\B@0FVQ>]ZdJ6JUbP?9LK,5HePTL8&ebCQM1(dff0,U>I3H@Q&?c1F3QJX6&<=]
8S/-M>#P+Q64_0]7JN=O\0YD0I>#[cX.\OXA>RGA;e7S^4)8;)B(E_=DRMFdLfHa
_5(,Q5dU7a4A(06cWH#VOW<++D#\gL32gQ_,PD_&]KF)gOOCPPcMM:fUR-XEJ6N4
:=aL\G4O>[6<U96[L/bQe>)XTYNA8_)S8E/V6B4O<)ZD>O[,;TJN6+T<U6[/gDaY
^O]@Wf+OP@:KM0T.@^cBbYb)8GU#HJ(V[SF8YIAW#U[R\&/CT5J(C(90DYVT>>9b
W,4KN9#4_V58CVL59Jb7DM_[,Z=7;L/OTb9:(2MfKbYJ6e=LX(^VO[F@-515Y3XP
V1N:]_=F+[D]bS6AeF^Z0=SJ-PQ(VE2-I8U@^?-GQC(F8Xg>4K<bFFBHeJKG^eLW
KJU8E0R,4^&7+S=^>DaEP-SYaOVHG&P_EY&KDOdH3X/MCNT[3-aCf<BW4b2>0^]8
#]?Y/T08HE+/XBM9J]+;:e3\VP,>HR:W>gbML6H,G)HP)0</-cA8cbVcFP8VVXc\
W]HSE0F9GgQVOUb-6V=2g/,D92Q)7_GfL[6A76&D&M#=,Ld6:IWOcb>=N==;MT.,
_MM;F9M4&-<_-8I/A)AK#1\.OT\OD+DWCS4S#]Me\AH_A2<?P#DC?/ZXdX_LL?Fa
G:#S\IL^#g)VY3M2.3)b3b&?QeY&e#+dSQe5@da(-g<;=&SIeEJOY;V2>[5#cb[4
-]Z5U1>[ZH=K@33OICGOSf158Jc46TEWKGc^/gKa=;6=67R>(5LEe7\?\g\,5R[d
M=7&6.UU64/_S3<2=<T7D_#41OZ.&O\Y7B&U+f9Uf[4>^#cW;&:I)R6JNCgWABQA
X-O#;A8c,-->gf\HS.f\6MY,Md3]aO^=GJ^?5M?9)gZYB/a9Oc8(=+_V.D83(U7P
(:@+0ZR)be^LdH5eRZ(#\)I5cX(Y?K_N#5.]FIFbV@E+g>>Pcf>:,dO+]B:B#_1[
Y#6M0:d_1H2;SH-U8M>]<Y6SQa]a<.ETVL_IYY#1A<0VAd.d>3N\/U/M]>/;S12;
Qe)Pd3SF1R^f,)6O,Da;12R[MLY^2Wg)=12/ESKZJG.TWG_:F7/(54,06+\0K/26
??-fXa0,fb-U(-/YRF?]->;[b.SgMdW)6&;5<@bJ8D;,&H,9Z][E3N.e[FO4,XO=
Z]O(,)ENK9egLM&[H;cOM]F88T(aKbV>->QH)M8U^AX7J?aTRH,8I^4:e&>WUP,)
XW>XV^33cQY>=[SOg&GO@AX/2f(:6A[2<_-FIN:VKa.eF5@fI@=QB0_L.dA26>SX
:QQ7=C3W7.V2YRT>3+W6d#;-[TF?.]V#IQL,ZKC:LeD55Q?0;B)]AB/EUBP_-]G9
D9>ebJ#]1caf4c00NE)E6JSe^1(&LaO5OB/R=b?1A&9I,HfG]3bHPM)Q?->6b]NL
Y.>a99W:/HZM_WLIELHg\>EOFFK=OK=7S&F(CXeISL+7K[Z7+PPW<KFDC0dI1V/;
aU48@HDPKK_Z@?A)(2=Ve^@^8cHS0>XKNgD.:cc&Ld#GF,+dV3FQU^7.V)2#g5Q[
B;GA(b+;F@.0[a43^U=1TF,UMaB11>\+D=&TaZ/)8DfQ(_7B>6eUC.Kdd,@PASPX
gIR<cLfJ([VQ&])19[S@=(T?P:^dLJ\Z/-=#L\VF=0KXcD[=<B@64).T-E[SAe;Y
YR6IE?NN.&<P27>EK3;;VF.+Lbd//cQ:c1)]ddJB05\,gbDNfM\WAa/<6EV:\cc;
Q;\S,GBc2>,4L4/;62+c^#@7Z:W@ScN]98WPS9WNC[.2[:d(/(gaKGd#J/M\P5fR
QA7/=gW0eA\+[E8ZLK&0ICdW/Y16E0U=b4\8#QW8/RgBc],.Z2[/FN6Ag;KYWN;F
ZeUb/dS/K4EA8+g[b93VVZgM9^2bB&<BZ>f\b,KRR@b;J@B/M1ZSTUFCf5c-WeDd
FWO-)?#-cIcC.N:.@cW.@2YB^EPReU>GacUCLG#^f\Sa2R&J4RKAR5GdUG&?F0RC
5V..bUTJOD/OH8F2_C^1R3RI=__\JP783NC_a]AY75CQdT\Z4[\b60W=BZNMf7,<
9\(XAZ[5H;=B9P<WB+BPbPVO9(=9L+d9V_]Q_LHEa<[C3&F>KKE-3)4#O@E4T_7U
BUAH)b<^L.RH)&S+34K2^;&F[OS6S^9\eD190B;+L7MNH\V>.0;LYNA:9\Gd4ZTb
=2(F3)FWTH5^SV&R,_)60Q@@RHc-(#95(#+/DLN+RFa:Ed?^6a&Be[WA,@(SY1Zf
CGbLG2@_MJaCBA6SJ&B0dK&+N]<#(=14a<[LFULTVGNYLD28,T:83VY)YJc6Cae<
76F/U4K_FJVY1b,:LZ1=P]W2a5S-Q\./LR)8[F6/>-PSDOEGE/42>ce_R6]dVf9<
[OGXKC93&JV/FUfaPT4@[FffWV7e;9;MF<&4+QXU,>6Wc5@ASfSJc7HUF6Q(;95F
gN&I#ZTRD82We2O[88H>,CZ^CHT@:.GHDOGE.9\gYU\T6-a#L&8=e046EDCHZd^9
MMcf>H\=gWUZcBLgUcCgJGU?<.IA3O3&;V<.M,eLg0FEU:39H:KJ,26Yg;--:aWG
=58Ed\(3:@0N44VAS&MZ5Y^RN&:6dEDacb-3B/a\REce1a/A.eHT(/<TNTJ@g-Cf
2Pa0>CW]Y+I+)FH;81NS;K\^,>IB297E4AEdeVG?H,&\>ZW+3?KT#@AU+INd;?W6
b.=.QU/8YEJ3BZ:g/SWCV05-#3ZV<aEMFUF2[H7\W;6C^F,D:Q7VV@BVdU.ZB_G4
D<;,,/f)68^NCE]THQH\_-]HTJD.,#GJ+B32G-JQ:)8bC3?RaKYGT>V_EG,XN3+H
OR^9)>:(928+Ac<EIF.#TK<Z6>-7>SM\ZAAQUA4I(&6Of86[/H<=15B/C[-]F@PC
Qb0TP;;GPBD8J\28?CH;56J\[OE;EE(U.,(O&.VYf]#PKSC7H+:73Ea-_cH<2gOT
cVO,@RBbD/U&^RfU9,EQ=Qc)B,<O\aPGg6/H/eKaN3A#,GgT&]5d-CaK4HQLWbF(
NVP?GZ0ZQY-E7M^O)d.;@<K&ULHUN<CM(@&W<>4]<Q_M<,C?@ZN^VDgMU??]\;5[
gf&_=R,]ega88XE=fV7,Hgb;bM^6<U3fKDQN;[gMVIBUG]7+VQKME272e9@_L@-F
_X1H4)O3&6ObU?B\LgdUPV-/&@?WO:+56\?,E?SP+>HAMRg\LFF@3=,DVdeO+JX[
/-QSG.;(_88F(FEKF7Z_[;]f0->aZ1[C:A/f?<bFf;_6;[NY\/7-MR7GG3I]7O;D
6(@aS-a6K,0_F#,C\#K#b7+)c/MgXa^Z.1G=28CEJH7I\Q4^M=XM;04dJ9_:^[a4
Z#R^e_#/WY^RJIgE?][9PAVS-=De9HYJMZ?>:BXX:M?]bNASI&H2FH97K/JKFRH(
?_@0JF.=8O8;9A@6a1gE^XLBXHLNQKQ8LWQgHf_:8JTG#&5DOEOA5Od@,bJ\.=N&
ZI2G@cJ\SVSYH-Y5]ddR=]4Yg.]Z7d\,6B2@A^8?fM)e\N@@:LX>K_a=RL?I&a4/
4F^XT,#\3f?WIBDV=5H54L^BT5<,+R<.c2)&UIaF.eUJb?R7.LV#:/UV9K41FaX3
S\,/</95S6dCdW5?P=d<^)T6I^3;XV\[TN.f1A?20PF7\/9DfE)/=\F[^?POfdI\
;d+J5PMQAK4(S53Qd.KGL[fb5;X0VK4JQ.,.6EZfE_SOeHOa4SY:3aJ3V-0b89YC
DGA@0QAV2E1AB01,OR&ZQWCQXaTK:,(eN<QPKKT8W:]UB-IJdB@gV2F<Y\&e4SE]
P.YHGISB5AVWg3ZWPgQb2bU>IK)YU]bJ,B)SaJA\OWPcI+JP>B9ML@)7MdXM6?-C
53_&W04Y_V/87X.P:TH6F=-3D\_]+=6cIYWFUd<IQ+?VW,?5=J:.KX(P?)6JLYY4
\3B34]),D[.SPJfO_@]@\,<aD0.M1.S7<S9:_=R+bb10KPaKAUS-.RA8Ud.K7?K_
]LHVDF2B<Wae>C7GJ-KQRF-5e_WL+A>M4gJ;K^_&&X)W^YDF1TO5F@UYS#21?;;F
e@M-WL]NW1I:WR7TVfG/<5/UQK>4HL:@.9M7aZKHT6c\SY29cfa>_7JB9#aVIHCP
_:<FN2<7QVHUeb(\a;>cC7X[+)<R6/8D6Z2=f(bVC818@Q^6\e\KT)-JN5[aL^[_
/^3&TgZ)P.M.]g@<C:bS#^9-2+G;Wf.T<[D&.L6/++cBZ^D#C3D5I:42PC:ST8_J
b_?a.K3F<9?_bXE,2,0-Q,=VP,dV60dUfdZ)7g(A21NXFD6W6aFLF+9W4+H?.-dc
9VCP/YV8O#0R=NI.2KBeLIf)>\>?8#K:ZM3^/1+O(@0Z[4@Y\C+KFfF10Kb7a^E0
::HMPY6<;</9YB[ZGIa.9;LOEFeTLEI-fZK3G=B7<Ba)49,8;OC,_]cQQf5)DJ,A
]T0U,G<@F\dSa_XT8FR(=>Z52;cd=e4Z?:S+QNQK?(YbOA?BP4#YL^^DAHDCZ.FL
J4[80T7?b=C?,A\d#Q[//JG^IK#\N<XVJVK+VF]D49V]Y-Y4ZFQ-F@3I44FHNCT#
?_HYa\5:-<D/DL0NLQ#La]>[bQK)aCHCQIW2&-CBZ12VOZLG05VCWB,Rb0c5bU?R
g:IgdT\+\U2Z=84g178O4E8?;&aL+?eI340dLB?CUeU:S/52;_gG,H]<[R:,eScH
&.I?g4H<VML8Y)2PbZ@Ba]ZW6eS7bT,&MR_)J^^G@&P\2Zd23BIe@G\[Y#+VK1?&
<SZfXVNM]U0B,O]K#\R&GcZW:=KC8gY,]82K\4@56B,(#6f5B_&_:c;JT2YC4?bT
)VHLaUT@IbBIB<&UMYgQg5Ob@a\CB-Ba>(,)OD5I)PYJH=YDF.ga6:Kc-:F\@-KP
F9TcJ\>^f:N/;X)&eZYYecL7L(a\]+S@BO,@;F:RJON9M\?YG?UXbe<=B(-I_4NJ
^Fb;=>8/Z<5gZ)DLEG_KQ>AI3ONReB6]\9(I9K-7<V5a8H85LEJ#/FK#/1J1(E[c
I^=/9RY6M2L)RUW/\PJ+YZ[B\U^GBRQ@VRIRY<O0]YO[M.YNQ0>?1Q:\;?R9#QRN
a5d97CS:g3?)SQ=)[@g8agb+<L8&R\]d]6V4dY+fJ8T88Q7DN^aOL9H+SB3TaJ&/
bUP\S0V#/G[OHG=)R/Z\+)04afP^f-TA9F7,..58-5Bc]X=FF]K=&>YO70XFf2;H
f4J5D?DN89?TXf>+UB[R&D)J,2:]\9BAH]?_6@C^DedQ^g6FQa>F=3)O>P9GRL42
A6F#WD.4;2H2S9?>57?A=D(&&R^WcLEJWb;e\#QF3-H+f\Cc3FeS1aA(_c<+P\>E
/Q8gXD#19=7,Eb=-7,N-QIK01:>1YL&S(\g\IO8ISE^:2aM0D4^R4[Yb>EJDRbe1
C5&FKPC\-\]g1=>S=:3WO4F6cgU48DT(f_K6GPJ?B][S7RNVCICBEUE.J;=4+P(O
]E-P>d\e=X,@88.aX0P:H9T.=[deLeG:@59IV5AggPE]RBJIB4EMOZ=A=JUX=:Y1
MJf(EB80&><@I1HD@7T2I\bRd#BA4dNB_:CDY\f/\#Nf4@;db8\LOWOW\Af7Vca:
0B6d3\&b^aXDU:=6^g#EeN6ScAYR)LeAG-Kbd#U>8/M/3A(\9gJ3^Hac/@\Sd7G&
RKeSD7_SGA#<>9eYPKY&ASP_UL18ACeC6==YAB>3Zg-+b[_1P,Fg&XfCGIF0[L^Z
>abTg#C9X4bK@+:,D.YXI<^K@O6=?DDE>Vac)Jed9HOa5,RXEC@8XO+>aK0N&Z9]
8XR:H0=3PLO#F)\?09DN:P0HR89V6c)_QKYVJYQ+#^AKIY55(.,;)gJPQ&][EJT+
>2M6@3e5W?AD#D2McUeK0>#MA5XbQH6>=CG@<VEI/4R7I(4HEU\FV(&-NE)a.Y^-
_V)^7.Z4fW11KC6V/Z6B]Y<F&_.4)bX]\7&0YR<?2XRFI[?65(>@\K:#YJ<WW@3P
C-RIfCU>IL@C4<Z)DZV=<P&IJW@VA9[VM-Mf6I)fD]1=eX:H41HM\EYR[bVI/V5T
B,XDaLc+O\/G0>LV87BeeHH761=9eW+@=R[.K.QO:Aa;Xff^YR1]:PI+3fC5F5^6
8c(a(@;Q#?^(<(a,_<b#.K4:YGeX/\91NH\]\/VJQ[<8SIGHTG.25-\AHPW5BBO2
VDU&17R>I9B0WcbfJC=^<\=OCKTge0Y66g6Y+)GWZG(bA:,WV7(_[?.,SL&ee;SF
39g\e@P(O:9WNT^T8Y:5JFCaH>If:1YV111Y^FJ=+QY/\(bRYY>PK53-B[<X@[1W
81IA<1c;1E9P077bdT8PaN_O01D(A2Y8BL8FZL)d)E;4V8c/P005]FJ03P]-+<c\
0Ifb3U9[O;J)ebK+Hg:6,c7dK1Y/JRMaC[7()C#ZKEL[\@#_T#UI2=c2^?XDK\Ke
/gZTQ/7_H92Z/L:_0:Y<cR)5+a&>SYg>Z)0]O8?7EK2C(@8H07.5?DOGEG9W4ZG3
E&:cS0THQ?Z)M.=f-?(QO1@MFGP8U;I6?.F][)A_AAcW.:NKBXeJ]^P<;3[&X)1^
5,]U-;42#,G>G0b>[Qg0e+<E2D[?YV-EW0,Q\31&E.-3PMM#ESdRFFS-_PIQT9Ld
S)/?g_+O^cBF<;#>WCXb=9>&3>S4:9.[OY1d,@NL+:C.\P5.S=@NRY,<Vb96ebD.
\J_c8>3@#FF3+6Od/M-#V;HCW=P-U-2F(8X7g,(U/WV+TRF>TI00OL+Y1BM.14-7
SZC66LL(1/g@@M&?F,VFe^9,\KIJJ^:PG1JM#@[2YMY2YJSR3)QB-S5S()LI=&Za
LgNf^7VF[,QV-M=QP[\YBY2cP10WXVXEFDV2V0PJ^1QM2cOS^<>X=9OU[Z,201>R
]XRK8H+6E-V8O5HU[K:\04CE20>WW-^W-0.@@8P[eDO0JQbGG@H-[X\GD14+RC3F
X&cA4-_IN2VBIO/9)/:B=[,4^GWM7?0WX,<]#F8#)-:b^UZPB5OK8eHN#@TTJ?d(
Q9ObIf[3YfUe0CZ<5/U0/A1F>f@+74::#9.<08>AVT@J-:#.f;6[^P:JW3D66TI=
(=ZM#g,]:2OcV<7?HaC[6FF^LS_VJdRW(gOU4G-SOf&P_,c2D-eJ:UI&OP9\L#P&
2L,B?P(T).\#-W^JOL\T_+=V/TCWC.AI2^624-f=Og;1_Ld(R8@S.B\6DcBYL(aF
ULHKT6>D:D.\]POf_,>M4)FGRX\0e7aPBAXa<c<Ba@XIE,+-/TB:A<^Rfed:-QXF
c(Y+>C\Z#W9DPd,G?gcR<?CA#A<)]OdS>NL3a:#O)Ke6_M:Q0-:M9/B5.4<SRI:?
@6M2A57bb_U]9XL:0+1@)/AW)f[#DCR^d>44Jfg1RS80G=XcTB7MWePMU&FcSF)V
(7BOYRe,&LB(\a#b#EdR.OEQd@2B[1aJZ)0;GX43_P+ONe)]3(.:B=gJ0g3O@DK5
fXaN9c=-<=KD3(]\2+Ug(5O9+Lf7<R-Z8&)/5#+QCFZ>SE1gHS)4SVaW[)cDLT+4
>,>,Y95dP3ZH&Q>#1RH1^[YF5>R<W][R?7_F1;M1<8/?f-OX[SQZX#87c(R&#@?>
[Z)2d;-,Ofa=M^JLOFOPO1d<)CW8G_Xgab2+Z5&+]a78LWdcH._9>03-(BZXSN]J
C_>&,@5S61LY+0H/YCe:Q9a^_9R3.]\+WWLE3\?DW&)LK\944d7fYUCX3<^>GO8M
V)+NWQc0JKMb<:<?_/ZS@a)EO:6G@]?I2PT(:XF1/[2AK[^a9N-8SUY9IQ]#O(Z4
U@gV[-\5d5Sf>AS@PD1SIbcH]<.a9XMZ-]8[?_ZTGU<fKK#JW[b(<K2I@BH#FS/c
<TZ)K@[.DZWF\e\USaM>@RaP@SS^0bGN<2,X,+f9UgLG/^#M+)Kg4MS3IaZ:EXY.
WH4d=W?K&1#ScWO-Z(ff&@+G(6Y9A^10EIVKWNME)]#>1N(@/GN)4:(0gc+CSfM>
I5F\^&<TE;+[CRDY:TI/](b5\Yd#L#&SeVIN](MfdZ++b9GT5b(/O][0[0MKHP/:
)#<:Y+>HU5D#_?G9X:W)K&KL#H&-HFeRcHQ7(\7T+K3?^DFB87UJV18KIcJ?U(&2
/1DCQ(WP@C&F)P?HNEfQDb#AgY,(a/8\Hbb\KQI0Z,K,KDfH7ZEGg?.NX11dO<3H
HZ__D?SafER1O:YeD8B:)]1X1@[<L4/?@XBWeAZ?][Vge9F9KZ8P3STILPK/BN2;
b+V#2SfceG#e?KaTCO\K441E;XRYLJ.f)VUKGe_d1&3=G1H7Y/.T3Q/R^;Be<=4;
SC24)C+g6#?LW)(DKYY0OI;cDL\M=?XUKFZ:<:W[OLG#6GC1&+VI=G>Qa8+fD+L(
J>DG-SSMOONBBPOg\AMTc=DKd7SdVcHN_BR+]5.AV][M7U9T2^[TKMKKCB[.C0c.
TL8a#26RR=N4>W9.[4\@Ld>g,W[+6d#&90R)dKFP0f/OU@3B-c3V9DDFK<J(?V.R
_CI^J8a.+AJ&M/9/JDJ@McN&0/ZSR>7A2HP_V-GddP:WO5IT8>4MG)7OfW08CT:H
GbJ+WDO>cYHfa]<=<TN,G4Rb.AaO4S+cA^DNF<V9fTP)Nb[)09PV&RcH0fR+QN(Y
?Y7ZG?De))_)2Ib63690#522FNL5X(_]e9M2J4#<66++Ve?MQc[dGVNNLR_3Z-4R
PPR&2,e\7:8?4?,TPZ.&TWT\#XFG3F7BR;H;)Y6e;AE\fOXWX7HVXXKaUA,A0?bQ
SN3:/ccWW1\-<gObT[+XBM>DIOB^=2TUAKf)05FAb?EWagf_8b+gd?SaW<AD@[01
5-(7?5W2RR2Ca\dLU[6PF4QJ+dg2f?I=T>EXHe2UG8>9Fb)+NW1Hb=MDS-g(;P(]
H\PD+)UaJ80#_BES-LdZ_<B,WZ]YIY:-)LT4F^D@eB:&YE9SL<MZVgQUEG7Ig9HM
G#U28d8((AB#OO3aP6DX)H]7?beOJX7_@TYCCCNe1(27[_/BVGO.#F4+8OEV<M>a
P]YgQKDe:Y()L89]F8^B,H&59J^f0Yfd\5f,+-KD72>A/dA7.a-.[1>BFc,L6DYM
d\[N)8YRY<<+PHC\Z+/AFMCYZPFH,E,)K].eBDH1Z26>2R#IY=AN[85>U7)QWSB,
T)N[;:IPbT2f.IV9+bZgWeJa6fM#\cgTN2F3;#VBQ[R18Y?1FH7X31,.4(PI5BOI
T4WW/+T=(+AJ<JZT3YIS\1744T@B@C;?\>M(DE/3gRC>]a;_aJW)U3^Z&D-P#SN:
ZU1Ka)]YT-.dO/<aOLgRF82J#/6g^<<(aHCH8I]g0<;JM[c]^OXG;;faN14_cZ^Q
7e2S6QJ5g7QdH/OL,3MY__OZ747RTL0SLNe3([9Q&/\G/XUKY[1\\2VO[aD\XR)H
]48</1HI,J91f2GG9/WPIb=D[B\4ZJYQE-7c;1N+M[MfY^;>^&#c[KX_+L7bCG)=
1/#J\&.=KBM-G.&)edJIXO64b2Pa5M;@a_/d34;>N@0c&5-MCB24N=@YWX<<S4<]
<c.bD&@@)<RLF(S>H@<3[e[9NYHXfcWZ9NUIXb.AKJ=V,DYZUf8:#+cUO>ML##Ug
44#NeOGK@N-DNDYZ.J+.1W^BHE-B>+#K.9=J]=\14S7_T:E)1fCbbGR6_\\7I+E2
c060]SB.0B.>UDK84OG[_EOD_?3AF^,5:&&b4_ED+[Pe7Q0e&S7@gT+HK#?3,LQD
(O#IWH3K#Rg?HT,&]?LQS:,M216c<SAJR8U?N:#?VeN6gN1K/X\a,;bMK;+:(YgN
8gL7H1fdHQ,7N;FX-QV2V9IfT9XX_6@TT8_F;?/,Ob[2<8M5^WE)T@EFC?/+]F)N
S6Xbd7\;BaCVgeBN^>.8+D9XUf,J(N_^R8;65-,C6)+S_CP0Rc5G7))R4g^1,W>O
LA:,TJa3G/,B&2JDcODZ:(JU8?R?XS4:c6B>\JN;+FRK#eWP5b#/MH/+3F+J.[4&
OL]fX0A5\^;6ZMSCOY(43V+f#G>HdGYfU8#>6C8Ne:>fM#J\gN]L:(YdVUO7KI)2
H1C],U;OZ\IM#.MVc>F\RNQ_Q?G5>58>]K<HAC-&\\<#=LI2]b>62YA?IUS\8gMO
K7d_=.F2.^D3M#eN0\+0b<Vg=;1POLH[g=,0&W7^aZVN?9NRZRNR7]/)W+Id,]aK
?C__Q@R;])Yf_FYN&3,LaL5,@#<(+2C?73S;J]X8AKN.af8\1CEO9^XL_CJMYVN@
6cWXQ<P5f1R_.=OTFUfPcBK7NU,^M]6/VQZ2fUZ[I#BB>]\)(9I9WDfEJ7+ZcN2<
ESOcDc?IOEY_2FeVE([[QU)X8b\bRaA:J^H&UB1[ZWe#d3(WTfGSU?(S&7G(>\J4
RM0P7<1<\F8+L[&E@Pf0[FW1D<0+4X]/g5-OAT5Q+Qg9T<Fd\\9WJ?cfX75,RO94
7H9ZQYfQ,2_1FO6?[C/V3=4;,VE^K\<))8+OIWYOLX.&&..5O+Z:Eg^H?Q-+:.4I
1@)MK[/\Df)LDFeeHaK<;=38+-UI_0&d@G&dL\+K+f8f)RZ_K\]?-\.CP0)6U9I0
\&UP#a5INd2f[N_51<:.Y9Z0\E>R-\,52SKaC+UUDPDTTcZN,:225&7<FNEBWX84
G8]R^7.bCUT#16O/[02(gcSg>COR(^C1UKM/SKQ\d38,WWK.,0\P4[1N:8\GJGeX
d5[(@dKQg[cJNRFVc(a]:@Sg.6LAF@R/c,X@KeBGJ.b2@,<_a=5ZfKKET+A#20--
eI9KBE^@ODTaTKTZXL:,0=a\]eCH5be(F2&XYTXd1@68B[>#D(J.cMf\<W>D#gDW
Q@@ES]Gd1KULJB0PBZL,SdSQLQ\e7AS>BFRK[A+IBWXBBJb[^B6?@9,XKGDG<LV9
?)cY1,;BSXfFZ9).<I,+_Je5MagS51dWfDTaFP4(OYSe6ge2_QgPQROc<]M2ZC^0
.F@d;>?MK;gRE&4QB^T.BRS=RA,b+ecK9P:V[NJf:47Y@67EQ&TgeLK7S]T92Z^\
UP^WOIMF_/S:-,^GO+f^.A?6Cc-KKV,c]94(G\=J)<1[Ic<L:96f7U/]_d(VP3JS
WXF1<;fc1:Jf]DQ)D^O0\=fa=,D:GK2PTN]Q&YPA)QG5fX)^RDaG:\(PZH3+@J:@
G+I,393]_[Cb;9JH[&^bfg77.CB5EE-&]?LV)](PE)^SKZM5Be<^D,)>^9#N^&&(
59<()A[G(C,XHXX1B_#1=Sc8;8)D[UBcESC7J>-4^[b+9gMP<A0.?A/c_;E6C[eV
Hde5D),B-bYW<^+6CKb\=Z?^I>;Y>g;3,RV:FJa4++HU7WK6dNDbDY[2aIb]4]]/
7O#M6556Y#Q>.[J<gH^R:)fQ1XJ>/,@GZ;:ILBT,G//CYPeBMU3fM.UYa0Gb12P#
-^4HN+Y>I9:.b_D.9OTW_#N.2(C#0A;^HQ#,8XAcQ<^fD<B[g0QR6F9O+)=XVN(c
:2&4OXC-d7=a&U/eWd(@]N8J>4X([>V?4?KP[TOUg52L<4D<,W,H,;BeXPbZ>H3a
D)=^DAbE:G1+,GRL/F[?XKd=]G#LFA(AXc)ZI+0JT69[.^E.MH7T?01#DAb9NCUM
]38/FEa)NRSQ#9=c)D\#Td#=TXaN2<R/3_cB)I;F2S1J.HI_9XW8J:FT-3]4+=Z3
-DT@FYWY,HV46FN6^W[+0-Z18?ePBLIA-=4XO8[-fO3SB(MgG^BgSWb/aE][[]]H
R9JC)7[5,bF^2@?PGRg#/^eJ)(1V?fW8N7INH-B8-.W<6cENF-18;M].S/216-O)
8PC5,]RUCL-\a?I0a0DL>PM2=-M;dWSGH=)^d4^-4[<6==8#FK;ZJXC11&J9X<LB
QZHW,,#b)N)b]NEWEZ)IMTV:+UW7Q#OaV.:,D&Y1Yb_M;K]H((HV_g^LL>54Mc^\
\J#+O:_P.)LD40fJ.[9f?=@7dMa(\A\_Gb\\L]F44#OE@3c_.7\2EeMeZMWX=JJ2
e1(1CY1f8a_NI>R<a-W]C<(]fageag,&=QS+G2,2;X+;A<g6Gg,NIBBU)D-\FW]B
?MCLg+7Y3?9/N25VX)RW,=:Jbg-5cbERE-@(3)AO08/M\/1K7+LA_EVM,Y0.&e)(
(a@3fU4>I6OVI9#<[?H/<@-;TEfM4W5V60>Z9G;O@#=5gRf1d]C&..V0SP7])gA/
Mf))&RH?@V<IIPa@@?D5&22YTO]]SePgG2-KgL=/?(K,3<1)85L0>TIa>PXD5BWY
J4X4[NdX4.W7,RZ,W>_)23e3L7_P.T/EF[[J@6U,?QG#(,F-H5E?/Aa&cPL?,9.8
Mg-;##IAe&[H50#^]>aC,:a?M2M]1b5]\-T]Q]?+C?;PJ<PG;b&Y8.?fY57-_fAH
G;:>:#JWQ-()70@fb>VF?VZM?[KLbQ#0B#GGG/)QT)+IJ8FU=dMAW[ZZ1Q(_PL+N
Y@9@^7aa^LU^/Y402Ud=:,4fMA261=F@:U+&6a?7+),^9/ZVXNd#-HE(2UI,A938
ae3(Z,UHS&9H;89NFL&MddH31/>N+1@.[8IY6:XT?YKYV2-]4>J&HdPdebTVO?[E
K/c.R-K3?5K3YU[5AR;GT4QXJ)7bU=bP9faHQ@B4B,[H@YQC+&UA8A/#bK1ADaJ2
2g3T[F;+/Q84DD3>F\=c&7WH0E0PJ1(fP2C-F)^FHR@+>f[U;M1Wdf1;dJ6-C/?-
;BWSfD:L/&YXGQE&E]dU<#Nc[W\71D8W3VOeSJfZRe>A-SH4K6KK[?EGFY(7,:9K
4J+5][b:S<6eH_<)<&+7)#F,Y\K>-5DI)K)+^Z@9U(BfYSCdA-\CC4I6?L/_#:^P
31,=VgHWH>:W.MK9DJ(F-eBR3-Pa,dP0Q9W7+_9d2cCGU8L3N4&O.:;g09J24L^,
N8c9I.2VKYJ&eTWeJ]Uc9Ga7^-7Qa.ERB#ERCSDF+(A#b?1J8UZ[0CVIQ9N_@S95
@](Fc=,SZ6a<C#KZ3^>,?cd(eP6b96UgGVg1O,]+D_2J8+aANP7Qf\+F2/]R)TLR
3S>+0(>IJH(Y+VTYRJ[cAPbQS)>0XJV8,8//b.SeP.LGNc(QP-D+]F2G7;A9Y>R7
PU&K53\bU6>H2N0c<RLcb>Y[a<W[0ac&IQN^JS^XTPW,P>GJ8/D=aDOP_W0M>7&a
a+@/1M-@@aZL-NUSbRASY(48a3SG+D>/OdJZ7bVQ(0We47L/?Y&T=(CMFKd7>+J(
2A1]c&(EFVfU[5;9GY7[-DRbJ4SIf3](EJA@(^4H?1SfY5Q7-PSDMLBfDK7DCV_N
6O-Q<K>-\E#,YA#0dZM93?#SZAdgO=)F.A=YA.:<NAXVR]+MUS?)UeOHd5CceU?5
,W6W@9:G>UMc\A\WegF5U(.HIa&)<J@A,2g,51[UGb4F#1VAGIEKS.]<4:gYAd\>
eUM3]_//EbX9DF__9]CZ7-QBN>N.dLfJW1eB8,)O30Y26=2NDJG1XZW+_XT4(YR\
903fdYg=;]?P+f_+HTPT-NI;U\Q:/JJG;QaA26=>S&P,5PI,0[FOS>NC9S+S9faX
8H5a3d8aZ5a3>?]Z]=D9MV\e12[eR/@0;OXZB,=--)8N=R/X]\T]^8#+&6C42^0B
gFB[F.LF^JbYCKX>?XGY#bA)HZL3]cA[/=V)#/WP.TW]Wb#@Qc@Q[GKLZNSW68[M
L@)/c2;H#?-O?W?5a.4f76QE5KG#bQD5-/I46@^TEIc1C]g]+PEB3Zg0\TND<_/L
_,6?5;XYP8N?0J,E2,7N?X-=-V#)_3JW.Ed2GY,<DY(2:>=&bD^We:\a(EV_JXcZ
-[.G;W?&6>]fVX?5dYIXOF2B[<=Ob8baGN;\XS?BGaO)ZG=eKS8D@YJ0K@)W3_CD
<N3.EV3@,0C#@I+^UNMc;2ebd3T.M?)OFP(S/TEOO#3SWY4/eL-\,??(2gb4LIV/
8QVPJXUf+GPGR<.44&6&.T:Z4ZeP9]d(E8QbXU<J:.aD3KU#&=W3g0+1g2(B8O3\
\AEbTg31NdS<5+IQ&CUVJ36S&9?0Q]=(eHH7CUeSeW[FZV>+4XdR-NA34MSH5Y[)
]VZ_H0N\A2cB(RcJ9P@1RBDM&TKIIOf3<&(APE8KAF=7AS)e[JG2+T4\#GbFS&[?
@d;2<_@Q(7@5TTE6cM,C>PKT6GUCL-.U5K&McO#4.9#D>If9:5f>97[16WKbI4dZ
7609BUEGBQP/Yd]3,MTY4[R96(cA3E3^-:2d+8g33:1P5e+AOE2&9g7)5V2W-PWX
8FEGS;d7;1NVgb9]]1E#]EeW08TWdNF#<9LNZNNXJ\Y9#\;_&O6f)R)-IWK(NCHW
/.?3&+4,3X(^9K]MB0UHa1]JRD>G<252UA64ARP+1WTE^@1N;RMg[cVeO>VYWF2[
VGbFOP>Qb;WL+6;[I;fR.DH:V@R>Z;LXDUgeLWPW&LM2U,<2fL[B4(-_7Y:[E&H.
]X(3E;IM&]U^G-_3f.G/M:L.X:&R+;V7-+(bS.XW4#2)?O/WJNPLcI[Q1FZN31K<
TX4g>eFPZG,bP?YPSC&7SO3gB2^+U&I0(E+UOXC7TUgc];5S7QGD5:A+PRAgZ@=D
7<X6PD<^MODEEV-&#FOaO&SD4D#HO/G=>IUZeEN1T6YdH,b90IbA3AH1C=46J/0^
SbN,1HSMeHdM/FIaSLMg1aJ:(TZ#4,g\WeNd\9a>W]\_N6,(]JT2ZAPK>=:SGX/=
(]7T.^ed599)LQ])\W(<6I=K7J?FF/D4E1.O-2SY^E<QSB[\V([^DUY:-FE@7d.6
gI3K;-5CY(3]3C8Z(aGWRaWOX<&]==4+;R9d7ZeceRSeANIPJ0TW<ES-57BL;:-+
fSgUB0<WCfOT?,d+A(H_P6A?A/ODX(S(;f2J-GPJbSZH?3(4Lb<NXQ+&TI>8S]0(
.&A[eAR3OE;_c=JMf4AXK#95[:R57IETEAHe=89c@>9YHP\9[G#;#=MfHPO6_2CW
VcL?QL,,g>1X2G7Zf#3(.OA\f^I0da+.W<5NW\Q4E5OO2DU7/?3=+=Z;JHJ<-Gd<
B1/]96FZ0MRD)fF-^]-ZW(g[82CFF7C]50@)1UbKQLN\@/ZKX^>Z[]aE5G3g9OKe
4W[JK18g;:8MT_aAcFV6g?53\F;[[RS_bCdU04JIMTE3R\Q&90+eJS;M@]d7\=Y/
I1ebPA(>.30/I2CP>SL@<6C)G-\L8RPS#T>0,YA7>>F0#Adc:GTYcMaBL:d]=<KM
=(O[f:7.?CYBKO-DcK2X_W,5HS3[)^TQD\UPCCU9fQ\3V1,g8@Cgd_M(aB^g_I#<
+GLR\OO2[A&b^22&Y.#3^C)S(QL1cU6d\e?W=<8G0H]XF4QM\3:db7FRD<MS:eOK
Z^[:[dA/49g)(e0^&X#W:^J2;&<<dG=e8e,Xe>EBJ4@[Q?J62KZY>Z^NHcWd91@L
(H>>#UTe>,DWgQX@6QK)=_]?d&96YQg\Q@)#=E70S<600.-NK0U/<6]:9C]MK(KJ
DRD72Vb,UO&9#;]CF_^=,=4B1V]WUH[dK>UeY:TIR6:L]HdTfdSL9Ag-8c44-A+3
geLN=]XYPQUN-c&^2]X=>>+ZJ)1@<g8,^Z4=:WaP7LA5e6^-&N#d<_QgXD2V(RD(
WZ[.(O2]?:L9Te^L.EC&-^4.Ig;&2&cW34<Db#f^/d#]RV^(Ja?bY38P,#JBc^K+
W#63DbZ27KGQL@)a8UP\@S8\[\;-QL[B-JD)6?YH)12Aa-09#83\=UX&>G>\Ebg;
/af_SQ?+\U;++7Na/bGQK0cc)eb6\_)@>\]FY8+C:e;=^2D@O-[6&2.JFXH3)c;H
J#Mb8R@&S8GIfD2^RB_>:.+0FTA[3Q;WV0=_J@>,ZZY-3]Q0_FK3C+][#@8#W/IV
e[<Dd^T_JTLA/dcAB/&-XSedG4Y3g@/HN]Y<S,74-FHdBBfYKfGJOAA0[#P.7((A
>:0DS&R[HW>6&aTS70@VIf4-EgfFOA-\Od;:/cV-3A\QQ30^K/_]PT8Y]3)gO1SZ
Ga4Z2[LQITa?:>5N&BS&9DH);;1[3SBKJ<eC7]]Md#_W+M]b_-WIIN2H0J3Ce8S;
B9,(,Igdd;.K3)R8#+-36NbPaI2=/:6JeBgA97G3LW?;aDLVOS>9BH]gWIWCcY^E
OO7N@/0]30W197K]4KgUN_,bIE)g-HVDM/K1L5]T+F[.JI&/dM3c_2W@?W7@/GIX
1]gQ=.1L1M@4c2E(M(/RF#6]:4_X-dFKfG0IcA/SF_[FYV8Lg]941S?8[DOCeNd2
f<cNO3QAQQ5/GG#O;(48&?bg2ONa<)]H,H[cHX=YD&44[c\18)-g,Oa?Z<bXKF#e
_<eLb)9g3fATa8H[-J](&Q;YG+AN+>JN9X2XXbaR)J03DPVI.cL0J[cTDJG./I5;
3,egROZ)VXFUE]XEeH84VT^9&\T_0V&9W3&-bIV<60EQe[;F.6H3>:\;F+S3CC/6
8EV\D<8ATE1)D.P4;:Gc\cdKLQNNBM\&,DB0-@:_:+L_a3>0/1A;/P1I^ceb)^GT
aI\Y7KYLeR::8/O4Q7_U5PXXU;S:VSFNDITLEWH;Y?MO4aQ/NA=F[eaY73ZgBQ3M
T/M]]F#=/XYQcE@>YEWQFST]NUY)69.(&8W8@1803VMQI93JE^&40JTYR0MZ/#g4
_OTOIM,;;b#IVS#afA-fYd?8f<LPQ4>AO=c+M9M[(/eW+<WWB8(0U#K9]V0=YJ\G
M7H^5<I_?V:^dVH78E:_2C#1>070I\a@I:D><42?ZF1NZ5ceZMW/=cbM\Y]g,JUA
=9(J1?0\Q7-D;#E:WNYQKFBa9YTWY++C;FFN>g^84CT27XLKN<E^TT_,G-5(_>fO
1T2;I2>WTN&#fE3=b,&8GK+=KCNBN#>;6UXCT7-TTK=7;E2.?QJK-4BF&>e51(U,
D+5)=25<XJ]eA:SR]UH/C:<I1bKS#TIVD5TW]88]]OYQ^E#/</)N;f4eR,,\7-eg
\a27V#1^c\\aZg-\/N#S5=fU9)GC3QRbYI9US#66S.W0AS=,V;88+5K32LMNgTEE
Mb78Z<6dP)5KQBX##]&6F@Q39>I-KS+fW:E4^4P=ANGcd&-<L^(3g7d7L+1#64Ja
K6YQ#6Hd?<)KF31Z(T0-cH=;RB)2&T+aO17b?=RG]<O]\3[f:E,C<5[5:C(@J<Tf
51^RXLQ.ZD=LgACSXW9[;Qc_8O@T7\:KRHFF<c>&,AfbJ8a,+M:;636[;B<Q>ARa
HC\8[?37=bCR?a+C&a07I==9YA#V)#\]Y9NNB1.LZ/cR/Y,URU(<\(K^e6b@3],e
/Y?R1f&8b.1JXT2gI8#8(GD\CBH;Y20gV02/LX#aJREKY,0(Rc_Lb&+K7;Z?=d)\
f.Qec\]IZO\dA/1.Xd9^MWB\e8IbSHK]ZPM\20-91]bQ@I@:6cOf];&OWaEeD#TQ
],]4)#PGY[:[.00C]P.O,L^\NXO9#=IO.X.Ig/abef>]4=f?b;5A<gbKOeWGTP^W
I(_g^,3QKW,1gKG2U<96:Fb/1N9E/]b-;[+9I51]43#F/M8,))]YCcVK[9bKPI1K
66F/:-eK/ZLQ/9EBfEJ:M,^IA3X9=._cP/85Y]K=B>+L;4+(aRV]FR?>C6MW-J6^
2DYN4a^UG#&cL[8fA?[4L/Zg6;\cX_X^>-JGQ6^J=B-3QgcW)\g;++1;Kc;&7WLJ
0BFL#^N;7S[I/H>V;^R]TZgYR&,fI0JPUW+VR>IMUM/S?L6EAW565b0D.HYE/[RB
3].R_.G69AVL?<c0V&>.1cQE+?Z5NeFXbU.DCV4;^c8F2KB4P58UeIU&)E?eHRe=
f:-K7f8cGM>M+G#J/HRe@0T+GgJ,d_bf[7^D3UJ\KVKM#^@gT@<LSZd#4S1)_0X:
>C0XHJcAO-S[B:bJ7Za+K^gbR6OOW^_1EfA6Y>38:+aDLH-bS\SN(N<Na?O)./5;
K5>Y^+@@YTZ(Se0/5aG\RG]Bd>+3A8-9-F=88aE\#;P<cL:G@GMM_7VcV?a3O,\P
A,/A2Qb.LZ09dZPT06agW-IWU\\G>=Q.YbI#&4O>-(#)5caTYU5YZaKP#(4]/;B;
4DA>9gJO[DZ]SR/9E#K<_U7Q\O#D,?S)2M2+5MH0e\#9-]bAO<]:^9>VUB]B(AGf
8:VeX<Qc>44>NC<_#OcX:V-Q1@=6d=@>IMQ;M@&A<0I](,P-2-UC@Bf9LY+-DEE[
?3RT3/.>O759cR7&75A[aD)Q8&+)2-8Y/CFf9a8?daPC/BTeQ>g@Vba_H?QfTWMO
D0g4W:O=98/:YO-&(-VTLXR-c.H:QGXR)\SJ>dW(fe;LA)ZGG#aU>c=ZNMDN-gG;
R#4e.>3NJAV5F(ER8f>OC9G<Q6de#Y6:3_FDE)GZI0dX#=\Z[2?gAY4B4T]9U(?A
dZIVJ=\/N)(e3c,8VQTGIX49#8<8)FB/f;f+V8C;Idb+T&:PR65SD^7;^QTTE-7&
PE1<_X<W9+:ZJ;+O@U?S\24;K?K>\ZPR+S4>bKSOU\==:IJ>d1bG&eA?aRFG9-M?
7JW,:660DN9-_M-G:B1YZAN?0e55#2+L7d]\99dCT<V&e87K_aLVN3#93NaV:VBU
b-N46?cNaGf<(]+3Q_I_\^=HP0a/EJ<X3?HBeQ[QPIe9D0a3TD\):CKHeJ>?)ET2
\X4P4<5&Ya8Oa<&9&=F/C\df01N+6MYU=->DY-Q-d?AD+I:cNO\/?@g[e/K7Sa)1
K3<OPXQV>TW,-C9YIWHb1Z_/O>-0EZ;dT3aFWM4;WEYB0S<:=K&__1<LFU)dA,bD
,PHYUb=NRFF_@7N(3W:5HD>5L(330>=]d(<K)Ie[DFL\Y3O394_;BF3_P4#b1d/.
S7AI3TGS]4&=R\^K<[9CVVPP8<,^>E1[^#3&/ff)&bI?OAZ3Dd=3Y1P2\T8]IQ:F
7T3@5g)UPGZfD)aS.0_<>3&.R33Y]UZP)^6HJcDCISQ4--D^^@BF_0J3F_8gJ7DI
PT_bCM;5S)X;RCNJO)]5^EV69WE;@#+6^CE@+\#2Y^@b6-_4D[57,TH,81LgQ\(W
5G-\4^T=1/dDAe-Z)#a(4ONM@RH0P^A<[W[U8/.AYYef72I>c_9)fMdHGJfDUJL5
=+<^c6Pd\4)FO+aT8^C8)7L9]5;STT#QB9V;BSCL5:EL&K5#(U.C(5F5(RI?(<JK
((e1c^\OPc7Y;BMT1_B,RCDW=PO[b4f0aK/O25<:^5LCa&aST+9SB28L\a#H.^.?
#G_ZHXCN/5;=(=g?V)S>ZJK-5eL8NN[MU^3eW3]NJF0Q3@cPLW-(]8KKO379LZJ?
-TE@8:gIaSVg2HFf=DRL2^b/EM\,6[AX0-8]QJeMDB/J#R+(\\:R=3DMJLgT;5>M
[IYCWba3VPbLD39ON95SA\_\fOBDWS25DX&I[QHUT3X+eC^98dP7:VGU+IOfOAg>
d)OL+L08J72T).;_^94XNP<@94Ke4AH+b0@=KXLeg-ON8.RH8S>?f]LZMAe06DXQ
#cL1/E[+[Be3@_aG<[_;WT(+R>U;].AL\;1B4CXCH[PBDE.@ZHc2(QF-HF6/7&I8
EEO:\,DY6R_FJR3N)M(^D.G,@,0f4R#]5S.]0?U=+Hc:;HHRfPF6+G)PDLT5<#]f
4fG8?bH2Fg<DVP+5<(1RJ5LfQO0]3e4U4EP3EM.<0-?WO?1.7IA]2EF)B?LN6V<^
A)Y6)eDR\V].1ES]7:[Y7_54JJ/Me1[C)S\385(+=55FWJ+BRFLH^N5B[]5Y8aFO
9?=<PYc(D]bU@fWX6\.(07PHMf8U#-M,ION,WfP5VHIKY/+[(DK<:WeY3_DQ]fAE
6-\Z7g7V3G+I);fO)bN57>]J>?MTMC&>\&8N.AP(cQ03bX8J?-Ga1gOTU2H([F:a
>.D3GGG8bQS]Q#?g_+L7c:98U4OVHDeM:O0:BT;gb_g4(2W5QbK>V)gY8/CTdD:B
V27da[OId)1;P3MUUSOFPCgT.4WX/U-BdS4O9E1Z-)2;SED0U?00(411GFY_/551
?E^Vf@>1E?VFX\9(cY=Y+<g4,3X(0<4FQYgGL35,0Re#If=20T,JHDQ_PdV2U^c3
aJK.FWBT7_#LNO,TGg<KT5A>6-bUZc&[(1035.K<]Ng]c2=HG/E5A.?H54QW;S>2
F7=>PW.@IM;\eKVe;,697GXagJ.K@6geR7fWT@VRA@])APW>,[eBb:T9U=gB\=[U
:8PeDB?K5@299cRE,N9F=S4A=1?2+g,GfL]6JG(-53BbF,P@+DV_f/e?.)T8IRKa
E^PU(d(4<0SK.<?U?GM(@U[6@G?IR,<edJEJ9C]C^\.\>CZ,@@4D;_\OHDT\dF]7
?5RNC=A0;L88+_NRTFM^:d.b,aFZRc^M-[GWOJV,V16&]OF=eO7;Eb3c7[6D6=:4
dME3MN>+^<_72EK/cL?0)0#JK9e4)?MCXZCA+/d>MYf164LJc_F(66#NY=eW_eI-
\2LdCY6BfFNe=\b<aF58]V=5gbQ@dW:SdSfc@J,NRP&7.Z-NP:IDUFO5+=[>>9e@
)]5G:WgO^&>SIOH;@d?64JH;f8dJ3.74PC6P[4Y6H.4(WaFU>^eFVN8/Y>G,KJbM
(ebMO<28Q9D)UV(g7@4\U,d_2T18<]5ZCMeLeEb8LGSe\?_V9c:PNW62Xa04[DS/
VCE]>8&Ea5F-+e/.4dD.3U(;/M.Lba_,806]VI&W@eZORZF9K#RUGe9@;a?-(]d9
AeB8Rg&TS(=128E=4J)FdG&V2JQ&6XM06\E&4Nb-0UGURKCP@><?;\Eb)_GE?@#;
I3.2N;d=X@&:MUa&[7#0#3DG/,3N:OK_/C4/_fNJ2HFMNA_UHM1=PP6f2AQaS,cG
]@e@[MH-=XY+I#IcF)LJIASV\+1IbV-V)H<]G+<ZV0/b.^C-6V\2ZJ:7.@6GO2S8
f@TO;N0eLMBLgMfcSVSJBXXWf@5R_:1L._N2>V.L,O=g62T:TC<XC3b4W[/)=L9a
RD?4HZ@J[5P^VTM9:#SPN#;T..UMY<G,([QX53B\LA>@A+^3=0@;d#5e,R5)Y5NK
0Q??bBX\RYYAJcWSbC\Q_WQ_9>S/7X.5H>e<e8Gf1YEb1Ia7_NY-9TWBBQcUS2Wc
.]U_Q+](]7]Q>9,8Y7/BL-a-H\G3LgL<E(>UTAF4PbgBO;,=:7<?,)Ya7Y>A_E)@
F@:aN8825c:D_9<^Z(F8Fg9771\1C1:^(^;9KB[R4OS)J?)D>,P5?3D5KZ)eAAM@
1.2QIZ;XGZHO4BW2M=_R;8GZb(8NEFTN@4)IR7.V#@P\[B@\:5:1:_eV#^/L09NA
D0^5@g1_#3KAcJ;aSNGOHP5Ye<VDgdMV.1Ue[.&>8gRSFP7Y]G;,;(X__:aLC.GP
g02^=8bCV^.87W.c:.K[;[E7(JYPg:+Y6eZ[IY;&\[eP6#C&D[&cT@+]6_R3g=d1
+WWOT#:LY<e,_-=S=<+V)]=0&D7g6A7AgQd0.M[QKR_PIDK;VP;7GBFPO?)+4-C/
L(77:10MQc;/a>I8GD(TD(VA:BLBR@)FdVS<2@:T1g._VC\89D--OO[4RV/^,@RP
f6dS3L^\A?W[-SPXYH8(NL_@;-DBgD#dD2^6)2?M,T4_JZ)#JfO3E()6+?>[VL6)
BJY7/&,(F\6L>7F.D-K@#&#+RFYXY&R]:3))U9.A=JP]@1L4C&,<]>b>5/aL5L7Y
8Q#0LIGGVfe3&SMH4-2McFO5?gEXNMZ8R)KL<[Dd/1Fc_Z@cP#W21GI_EDB[?U@^
dLeQ)RJ#&EHfVM8<:\Y6)(@<J3#K(GQ.X/K<PaVV+[d,eNG<PY.&BdO8<I,b+X/N
)YZ-FD>fL?,RROag#.7<9,=0HO#8ZLb0AVD1_3.bPZeRNGA9<-Y_4J?LCLHR>1XE
YMEOeMd:P&SKTRTLZaW?6HFHS^0@=;E[B[K=M3bU);[THO_G]^B7:DK]ME215_dZ
^gK?7C6,FKPXgN<5b-AFY31GE([\\565.X2+,1/\J:8TD]NQ@HI@2_CbFNU<5DN3
L&MCS1c@:U<bcd;R/L2#I+E20&X.>)LMR48(Id7Jc,SR\.D\;-CQG3_XQfZV_,U:
.MgF[[<>6K8gd]:a6K6O/Jf2[AS9IbV1c8W0a]9[Q_T(5Vb)_XB=RW-ZL^PB.O<^
fNQ=I;US35&/5EDAWf7dX_EOgZ83&@BTK&7Y8c373Q-Q-<f.gKV]63JJYHA)#:VP
f95+Fd0K<]P?7P8K,\L+8.WRQ_C<Ua[9,H^?UKISMgNHX)86/,W6R-dN+Te^:gV3
BbGYDE?@>O-:+a@D0:<Y[6JL85W/2[)A<FQOCLWA:/ZV]:4e:JPZaRAXVK]FE)ZQ
8gW)2b9DGO,4+?.W]4f8eVe=5(cfYeE]<I^6Z>)cAQWA331e;:-X-J)E^HbM_VMe
^#O7PQGUF_Q?^g19-]fS_Z;2C&[-a_4T\2fDUL/212I_G#S[2?VG_JVTB.CV\/,)
?G&^NQaaR6(B45N6ZZ#/=D^c0=+&fJ=+Y)&Jc9TeNEEYbg8gB1J1e<_1+P+_JW;7
44Ee_6Z7V2&DC[Q]bJcLA;VT5Cf9DaO@f0:-Z.:POY//^b4,d^/O&6QVOGMU6c)b
f8MGcb739M<cfGgA]P?7SUe9@,1Tf>bFS/?;Re=4C0.X&-&49(>dJ7@R.:9M\@F(
VPYSd(1UZ1LD<Xd/C>.g&86B0[4W4&_8(\MK66c->gc)B\M12:FYf<AB_4F=)10O
\,HTFRdQa@]GcO#Wg,H6&1B5>Y=)J-cE+;1J.@62T>NcIZR-BH=0O1E:]DCg+<#6
MJP_YB1D0TX0JM]4UJX;T2:f9DJ^LE_7?J-48[0XN@[.0J66\aN9dC,H9a6O@ZTM
9IVUN.gO[1MFKE-H<J[2+-Q:e(92=(ZAEVX[4cgNAF\=;=NI+<c)4JdQBe=K;NP8
Gd;/R?2FA[R/#GD#4+=AJQ<gb,:XbT.A[2&=M[+-)5RgMbaFbfH4YOWgEefc2<Q&
Y98K<BfH^2QXM,)?7CA[RR/gUT<V&\_,:[6PAIJHT@20.dHb\+L-[Gb0_aVA+;<&
dJ^/Ug>H2PLbADQBc(H/?@,E]JP(9H0.DF35GINQA_.@]>37WaT@YdSYOX5GW6B4
RA<;,(\M7B>5Qd.=(9__Kc/QL,XN<=\dS]2JZ^@-TAXMMEg91.;@#g(C<fYR:9C6
A]?[=H5)D^.IcgMW)@P>/Y]ZgA0b\_&[^H6@=E^6PcJJ5V,,IT=EY<VeRP=_MXUa
cJ>DaA]3+g1IX0DeQ_YXJ)Z@F.H;,M67/X[YbO^6).+dVFBC/>AK3X@=0\dLb8=K
0=)5SENK69>cY,G5?F[&2OYB==^EQ)X9#cgbeB<_RVbgLM0CHAZM)g,^6P=HVLW3
_F)Uf8R].e\fM6OY#73+DSgD;C,(,D+F>/eC[0Y567U@\.C6f2E65\.DO=1LP:TI
5SUFDA02=73Jaa;bd<_BS8-QY?4\dAL,YWeL=[f5OLL1M\#bR88U-I&C7K9-?@-F
..08F?5c7b,JRCdQSV]9\^>L_X;cJL4]QbU1O2Bad-gRFg\I)A,d&OEd9gfAUf-5
&<8DUJdeFD:JL(K1/ef=-\[3<_4[ec6.<:YNF.F=f^YCS-_g9^,R?C&?gY/c5E,1
3R_,TAV-;6</ZcRUNX0JD@NQ;gB[7=7YU<KZ&aaM1YUK,>Z5YA+(./+B31(Qb-0R
[+[WQe+Ge(IKOERQVdfI.J8-cD-NcTU)Y66Y/QX@;X0\gOd[;>Q)c>R=PJcb8+<Y
>E_YFU<4WWT:L_US?EDA5_@#b&TVD[M]Ca^<?-@@5Hc>gH\?Y#?8aLZe,4OYZPL\
OGYRXgWaVE6E(4Q&UA3<SaN6K&/1>/=>MP-I/I:3Z;0-4L7Tf:PO]cgN<P)g_&5O
PaCW24>#0>?XD:A+HQgC[a983I@(>8c@T#PZ]QYJZPc_c,fSfLHOWR#Q(:75+EbZ
HJ,VZRN(2E);K9KbeXU/53QCSA+#NFbX\/EEKIF1OIZB.R@ZC68FV<a[.dWUMQb,
>#AHPKa;YK:Z+QPLUfN0MZ[U)]O:-f&NKQ(TaZ>^&[1_U\I5Q48I8L71Y(cPMMSU
I]IU^:Ia>#4N^5OHgcVUTYUTC026NX5=7B3bc1(D9M-LTM@M,@7L(+Ce\E=3b/\d
[7E,Q4fI^O<,CZ^F1aO)Qg^1M\2R_U39NfMN]VPB7=9V,dB\dVV(XA5O;^>-:JT)
,/LR=3T9bIE18;=^G.FW2/HJDB/7f#FJ,5@aPMG18OMd4Q]S5(+=[c_=EUg0?>>#
.1Z2g:D#&(:)KTV3U-X\aEa:bR,+HB6aO2Af^&],;72,#(#B_W7T8U)Z<>KGMDC_
JPWVRRX.+gefa3B?-7]3E4bNNNB7NgPd5ZGJN:&7d(7;,D?(dD+e^HLXEDCHbB_\
GP[^9d0ZI<Q3E\<]SaM)1N4UF]184T^T.O:eJC_/=>901f]A72AcEQ;.13RZZ]7c
DM[+LfKD@C[,)[1<D5f0Sb@A/5b4.bLD17C6><UEd17N-P\e)EFXe5A//gSD]TPY
IBP.I?9H#7DJM9&GcM_fJ3a/_81A/T2Je(]]QJJEJL70,5;0X)Q>O807BFU_9L-4
U>,O>5P9M#aPM>.?8F?Z;+(?^^.&V>4A<E=N=5J;d-VgTRF>NDMVOVN34)(;5f7D
-FX/(CWX9<BT]@DBJ4W3d?DE1FAC_,CL>Q.ac?+,)dU>AYg\\SUb)8L1Y@MDQBQ=
2E-d.N/9cgM=:M2<EOeK\M3\b<Ac+B1SdS503AO0-0C_S26J#?DYV3A#2bRR8,9<
&e)_?O\WES?,[bDL]aTVW8Z(/EY.ZBD/Q#e<(YP?@AS33TT5OYVJYI+gFGC1.X:R
I2-3>dE?5,J)G>LZVC5T^.S0#8cFR)4I@Y5&NT:5/Ia>Q-3G]]=T<#X7CU7&DIBB
]RKeVREXFHf,VdS;W]WT7P55a3^]UCJZ_F#JY,-GP.9OC].IcXQ/eF\&6)U@:W9a
LF#_HR7fd,&N(Q4O5+LfHCW&PFL;@LKKDSa6L597P5\L[5Q5K5@]Q;SUT:QX>]g.
/[Y:H5A5Rbb.Ab?HMP-^Q0O;U>8VJUKPT+EY(>0F2_)OJ1GE-<Y#T7c1_DgT+CBB
BDN8PX)L7;9<N89;&OK/DQ17]f3.+1Ag:B=Ic73ZTU.DDB)gMUg=GOdS9e>fY(56
:JdA#b6A4[J&\\;PB4Q+(_7I\;5HGg1)O&dcUANC-EPH+,C5@NN5MGREL[c0gdEI
g(<_9CD/Ae3@#PO#CMI)7_VZDP.O2/JKJ(,CQVOP@fTb6K2AW[eag)(=FEKHYCWF
7>Q/:9+#MfVD3AR][Oef/dL?2R;WWBFd9MdIgBBC(I#Wa=DdS[UN8EAT5>=ccLPg
g/;E^4c/[6df]@?]>@BT@S;H0&8(;\T,#V-X_9,E2PbI:#0Q-]G@7Ae_.+PfKSUG
C^U8f0XK(LKD.?=e.^3cd^<CfV=6CRQWQdJK8ML-N4SWT+NaNUgX<A51I:T:TNb8
B)1GU:0DY,2,IVD\fK>+3<TEJb(7W<DA+6,\?:T5NY6dgJeU-6LW)\6EW&:?3]N6
F(W[5Bbb:7#\/7<48ZZBd-3S.^_E<f5fNU]TcT@([UQS/Q6\c:bU;4[(<D/CWT29
d7N+45S@522UcL[f49DcH6bf&G,YLf,W+BA<K2cH^SO/?8PfK@CLBaV=NW17=;M8
#.JOCY:^HMVBV<(3.Q(]&.@dV\X6<>:F&NGC2C:\@3P]_(&R&(#W76e828cPQ4]a
=9-U@_d]=)2UH&ITL<5J3/K(#__1QM;\Z^<U<Ga@(SNEVAEQEYWUL=NLK:S>P2+:
^f7VTcGG=LP7;1-7cA(EN)R(_fXIFQ_SbUE5CCT/GI=-0RN)\=Y0/)[MEM,dE>+S
K06[f22Z3_SOM[CX>[#UJa;Q7Z)bVFF_RCM7>TPG\;@C&A;3@:PR<D)F&RS\OTQ1
dLI2&\:4E@\ZM18F:B4=7GQ^8aIf?ND-b@K/M1W_N]]fR2fA))_&dQd\a(O&XC+I
58MDR\7A-F+0)Ha<>fWP:4aC22>\.-FYJ;/E=M6<@85[agLC5[TSS1ULDe,)3@/C
KVOWC[C^]ZK[-RG#=OH2,-BL#=I8LL,-1Pe.JaHN>^(FPN+5:E[GNPLa0(62Dg\c
9b@8\SeWCc[bC.CcS+)L,-#)/a#g/QWXf?7C\Q^Y0@OBIebK81d5?c&ga_RP-\ZN
^CHM:?ABWdV[T\f)6J?[Vd51#^\S9eO[9ZTbK8aB_GAKgZXF;?)]]ML.[3Xc,_8R
8<.#&?RaG)H<&==YHG8]0KF?0[V_&+V@W[F+2S)1=9JM<RMUaeRTQJY6SP2]&gA\
SOab&9Z47U9KF0PeF:Pb-b:8\R.[##M/d:7UWaV7_eSecV<>R9fO6H2(;;&AEP/^
aQ3?V?,@W7MS[S=B:eA\2IU.c6+Kg2FG)f]_)@J232:??7O7O/_J>K^=G2IaN;3V
05@?4X6PF-)85AAL^95E_c_\[8WHT]ecV865=J)15E\8Cg#A<(UAW7XU:GLNeXWV
2W?583MZEK]IgR(4.bEY&\W-4CS&D29-(g#]Bd?(_^D>;-.P&(9MI00\,R>.-U+F
c,TFBU+A<YPLR:4,fB>LXEY:K]Y9fJ3dWY/3L/bY_SP9UM(4?@ZPE,HT4QF;HIA7
HAC)G-c_@<T;.@]N11\7TILU\L6eV_EV,T=L)&b4Z09TF+3OCN/AccR>Kg0@_?IL
<H^<Kg:[HZ#V:)@9J^31U_gVCNAe5;X.:BR(b2d#2a0D;5C[b4?La.S;[[R&F^NH
UN]).^IbN/f_X>EbSL15&P5,GW_#6=f8^(<b/:<5f+PcIG<)2[XaKZf\@3E=N@8I
];Z<I]3\/MUMC+[MSOAU+P(?YGFd@RD?8=ggMM9ee9,gAWeGJ==F]-#U+d._P@FX
),4E1921+5MHH9N0[0DTU>8?1A2[F.+_DIG8#KH3d@.c(_gQGL9<^<LOTWVHc\/E
F_+K1LXdTIga_I>6R[S/Y(dR\K&0AIAKW18dO/T[-?6,3M^Z,A1//gcb8[O:V4K)
?_X4OTF-cOD\5&E=a_(VMLD:6))2GFO2Z:G87e2.fN_(:8F0_=A7^V,4Q)@VXU:D
.=]2GDOD@Q6I3/RZ6Y0&IO-+XeMLX;TB5Hg7O&QR:-)\7/IF^Q[;)#CbB?Bd7R7E
d68c2U[^/fGc/RXWR#RQ9G>6U0<2&J=Z6cZELCQ>=D=R3?]F-]Ta7dX)&\;^gccR
S)O6CbYKaDSH]DG2Ta?33,UDF&Z>O<F973:63f=N9/E6KXJX:-KRZ7GL=8F7&Xa9
de[-#WTPT8D)]92[V)SdP(PVB:.@dH@<L-2HZH#DZ0ZZc15g#]49EFP+0TY.]DNH
C5M2M=6.T(NI[3[@Md:;<d/6fTT4F>J@+J0<?g^;&#aJ.R[Q3FQbEG7]6MV3/=KK
;cW;_YTcIVfJ36FII.K.7JD522>89,<8HH@C#>?6UMb=9YVRMPI_F]a?+Y;CAD;G
((@P9AO[,)XK8RKLD);5YG6Ae+(GEeZ6+RGGC/IV,bO.D1O45T4U,<I#^Ga?Za?[
3T0:=2./?E]C#[B8IUITJ=:LTX#5HT_9D-_Da^;A@8beHG<^\E4T,T&_TD)UFDg=
+<;#3cBF8#SR23.PNN4]N4/CC-RUU(B>aePWbLDcTC(F/XE<&[Oc/QTUg?fEW7[R
.1O1>SAOMD/+2#=A(D:)D>gRd_TF2?TefGQ5&]M>Ha<.>7DI6814.,+d3X[g]LZ6
-HM3Xd]T5J1.^>EN<J?CG:301,496ba:OZ(Me2B&&7Z(YKC[feR<YIF-bdA+K9@5
@?XPH/[)UHa]K0:\6V5G1-FTRHWONK?+>V]^QT-.aY->6(bXUJE<[@<9,.1U.B<C
5#8L_^C[.RFFGH]MX3cV41J1&.f6GgUd_#5Z<1SC#Ve,gE]P+gc/KYJ19d\ZID6.
(<Z7;FeRL/97T3/Jd5_<VQB?]R:X800@#J:8:]-8BY)]0:&J=.DcPJY;9.IAA/_2
NJN5YP.B=<]e#:XSWcBdQ=fS;6Z=b>VBD7ERB=Q_fIK)U-:U9f4UOFG@30S859da
&#C_ZGD=?>Ve0RD&e-&2G4&3^<:cNTg[><@R8QFXX3g=@2QC&6;EId<fS7C_TC&M
3_L<^\gSO?IL[9Z<^61:dS_G4OTKbgK,Z2ZS_S7P:W1@[KH<:K>Q-ARR+3Q@L.aC
gbG-CD/2,WL5?0CJ+PWUYIb8bAK>A#[)4K(@V](cBfN2RHFQb82@C+V#4DB#SQ2]
LL-Kd4+2V/61#+bVI6B.N(Q=0L#.WMe06<1_=<BW,K24cPQ2A@+WgF8:SEN0S:M>
34,[KTH22?VdRdQK7C35@)5S4^.&<H3-XXfMaZT=MU#/M6JMB64GV&cdPMVN\d;I
Q?WE)3>a0ER7KY]YBXH8(P4O?#ScTU.7)4<ge#g.QbPVaD&\;S6<WT)/HSXKRF;C
QYEL7JW:PFT&?J.GG+XOHZ+G?>MA\B9VY[cUE8#(g=T_]LCCSdE>=LO?^gM1U>\/
_Hg(@#X1TW.(=L(;AL+@Z<IGJHDEg=/LDfAS:RI\aVWVe)CPbB,d;M;^DZ,g#JMQ
;d@R(AHUFT/1c^bBU&;^MSa6GfNdfH,H/__3LDB-ZR4X9c8LeX;ZeHb6f-N2HP1;
]3]c36]@Y.PJG6UH6Cg\+Y)NLfS/NJ9^?2f2fF[fS\^K0a/(LfCCc1OJ@[DA#XR+
Hef]4@IYZRXcOC6LXU&PQC0gR&PN?gZ4LAbLeeRaaM^^9TA@V<6KB.MdH=O,=+U5
EA&=UBW.^5B7KcELO.f0+MI&4[\W6X#L5Q&_93:5)4I>R&,c1B]ccF(4eX@dF>g)
UJ0<-5W-g^&LD>?S/-V2\.N<dARW=CU1cS8;2<GcB^ERA8<0FQ,BZ7>.AZ3:OMe(
PD0H55KHbWd\-G/aGUN7,XZ9PE:41Uf4L(&HC7QZ+WISg6CQ[Q4d1L#8Ha9Rc@-A
U4^Y1R^\>N-fa>Nf+b3\^T1&E2,QS<WM2Y\d+B2N<MbF4HeU_(8_<7EVX7>VU[S1
0<(PX49,F0Dc?F@X<R-;aQ_=L0-2/#]3+2JVU?CGQE94_ZNb\_?/O?E,V)5fSU;e
B-[DHDMO\f5dB-_?A1R6WY^fPWB#8fW];(SNL(_PWd3d5<,BUXIKZ#IM[@PYaG)M
HG&0Y5gQ.UBY9.W2cC/(4/R_e1G;_/Lf&g;&O)JVIL3(C,\XW_CO:2<\3ITC:2:6
;M\MadEO^8Z\H_VC5@RHMHe:V4G/@\X5PQG_HKU5SI,Y3.K4@UI1JF;Y>:2O:0ER
GB<Q^IdPHD_\YR22B?,)GgB,6+N>e]>QZT4#R_)5+-fG6#8VV?^Rc/79g-eD(1YL
GNd_&Z;fJ5VfX:Z+UU=e1-39MJ#@H?d+NM\?6^Pb=V@/[Wb[@LfT2UUH#+gYQN;W
QL(_A9>VCcY>K5#0YHP@IfZ,[>SA?1c,KYaLH9L=0[I#=M)P/cTcZ/G.CC)+D.HL
USKfAGa-)=E.OIe[CQKD)X4[(?K85J498FFW<MbKFYZ\;<NbO7@I-V[ca;Z-,Zf<
O9Z3bS758TL6cKO^JZH7>IRZDC]N/-\A28J0.>><1cR0G^&c&T:YOAa_[KbFT_=-
.U&86.T<YOOb.V]4]H=KEAZ_[af#H[S?+eWeX0:Q-XW\0RXL[YZ&;7(A;QKSZ4fY
AX?&^+)2[:;073(+&HPAC[Y&g5g.YQ#@.1Y95(/+_QCb4G+)\B+\#]]<O]7dSWJB
72F4,c)^+&P(IKSe^#\CE<=.F1D8L<K]\Z7R7D9U?d:3c]G_bZ2)3Xc88&I=IH7>
^?H@OQg,GMGXH6EXa;VNL(#A9T0feGeGFbd6gH#cE>V@4U6Z4\2/ZX9RU2LDQ]0@
ZU5-,O@X)KUd9#T0KJJVMST^8fR)@+OS:A8bADZ<JeVTG?6Tf6OD=)<@YHJ((S=Q
_(UD]Cd[AVI0]1-8RKQ(_>b#CNd=6cT1P2)QSbM9faTSK2+J2KN/fWJFfOJGCgT[
(NXDOZe\WaEA7^_bS=geSbgg5]OSe3S[M4KC5DQA6_<YF<_2MJU\\GGEbALF>X+8
ZYSQH:>;_EC?2D4TdN=<B2/4fY5-M<YGGfQQ^CW?9=5D-g#g?8P]VIINW;QAY.-a
6d7N:]RfgR=GFId[#._LF6^NB[I937Ye&+E>eM\?,S0c8N[[KNGY1g-,-CgS;^[B
bXHbeefJ59Ve_\7<]]b[N8,(T/[#1UebJcag+<QUeHZ=1+A/9=KgC7bCUV1gA[5W
G)3/.E;#eL=U.?89D2NV:bWfQ,S<O;dN)LUT#Igg?#JPV)OQ>b_-RG\gH-e95LH(
gB;)>,9_GOGN6Q=#Q3d7ZM1Q0T4-@H)Mb@gCPVZ=(fR08_\d-9<B1=5b^=QC(2>d
g@:6(JZ47W;TEfCO>\C=S^SDA8a\W[W/;]7;c:E50,#URJ_GC>V-+NH=8]3S3[Y0
2bWb^GV27,SOAN(&1BASGPYdB,<7WS(J.aFUEYaI1DHgR(-22O@ZZ>R8=5?-^XED
SFc[.V)KL3Y17FNK?ADR(&gHb\IA:J)35B#0F.O4_OC/cW4[S<80<L_&F]C0+85c
dVb6D@,>,6^CY_ZbI^R]L8C9agW.B7\;LSf6SH(NY_KQOU[</_36:&.KeCN^b8#0
<[./^:6@(cNP4]F?[MFc.1GL._&A4<8JgCKY(P>-O<f7H85\2Z9>G9bP[#A(<5WL
L@TOV=2ZcDPF:[KE7XM4VM4g]K?_887fT.2N+f<a\0Qb#9G7<7>.>@[gP)HX(W:I
I)P&X@&IJ6]T\7b1O.;?->@S>&5<Oa9Y+[:=2O0R:<6eQ)^I-\PfVKH#f[M0&Z):
?EIO#0A9:?#H)DP\4O:,=YC1G:H&+R(bCSK#cDT@g)3;/\NDD[a)WHB<)(g/D<H;
D\)P2D2(+2=-H3#0#e[#-\]Y8aOY?QJDVJ0V(4cc6),SX&ILb[_=7;^\,^9gBPQg
QMIRDQ(IDeE3B5H:F:8Q4g0>G7Z4S#^G9KY[V^IN8HLY5^Pa-PcYUL[S1,E2_?J<
,OaYcYHT0U#I<L<2/R^H3^P-(F=K6U;L7cZ.1URAEM,5/KaR=N6A&L5-MO);c9[0
1YA@b#:g<V\+2(.BHT<9cG5YNV]\\@Q<JL6,J^Ve>0^PJY1Z3.O]819g:U#A\#V_
\6WIX5V)acF.UJ8SKbL/OL1M[ebB2KeBd@3FP,gfV+[dKM=RdYYM55@-CJS<EQAJ
01^\)[)8-V-_3GXS[SWX?Qb7]OX.[66MCc_,9cNYE-DU]\fMFdPE_K1:gXA9)J/R
-)R4:Lba@U<,PB4UZN7B:P/KEMSNF:IV=]Td=7a)N6K-bg=fOIEA[e.Q<;>NB2QK
_&X=[f\S;(H>_<0\KT736Zf3ZX-/WU#YHF-KE1\R0:be.7?eB?IJc4GT]#(RUPLU
>UTFKDO]gP?b@e^c]N5+<FY5(Z/92T0MT_+,.J)J=:Jc?<Z&R7F7N,X/J83J;1e4
fWfTM987PL[,AP,+a430:ZJ,Se@-Kfb.7,AILbTc3Ag/E8F?2]M01=2CgLX9KRDQ
J^(I1P-dQd@dC4E_VSUPR8^MCN82764SLM@D=G\;@,+ZY_(3DXLfGA9-R:GS=VSE
5Y41e&d/NLc7X-6.E\+bS@3.,OQE?/HBd8JX15PI<#A[M+UFKd2Se,VbMB(CCCX)
bH4_U?B)0a+DSBP/<cB=[,fUIVX/W]QRYEV_b;_>/BA^,SV@OL)BdFY[T5]_2A57
YY,#aOE+-@Bag4;6M:Vf4+NHHQZKFcd\gK]6-.TP^S9/9>.O;:OQ(6Z2B<AROdBN
N</:<d;+aJTP6I3N3J&IH#2eT#F^eXCQAUD.4K4/OF-4a7DHcCX0F+1YaR;YFVN-
+YW[ZY[_#=NIHH:&K1IS<TCIZ)\4aS>Z,K6eGG#]eU2WCV9@2B?D@SFPQT>eNX+#
/Vg)..=])a&_>]FIB>=TOQe@:a>E4R^]515XPBI.E5PG(AS8L5SgHOI^1gT\LfB_
W#4N^:@Z?SK[34\40cVSg1>OPMQ^[>KZ=5^JBA;;SSRVLQbIbK1>1#:3?.Te<UG;
B1PPa,7&5UB[R=&gSKZVa/)P8C?8?aVGC+Ra12g.=]3U2@_K):5Y^S>:)62@RQ^1
<AO,4>L@&/g&@WY905bM,?f)F.#31;3PKdVH=NO@##B@V6.5dH?VK.^@3>F(\0K\
R21cb]IO1\L6Z]@H,@E&Sg38UJ9b;CZHGMAE9-SRK36E4.E6@<NOG;@.8>@\;6-@
/ab=L[Ofg(\W/cWLHaWW(<+XeZc33+8L][eS&Z[fW>&FW?YQ\b/A88;+M2\I2WA>
/7AG3EE<#)AdS-VBD&^VPSb9(8cG#,_J4,P,d=YVNQ3^D(5RdW#acJ>QH]\f6?VC
c4FD?>WFM?dOIEZVg@HVD;5^.-TWFL>E@5FeW&EXMfcT#S[ZQ-768,^(./P:FgZ(
,W.7cN/)H6&IR19,6-G0<&D4H9D0<S1[Tg()K23A\e2,CA^1g6A9BF8MKa6I[f/I
8&#7IM.RE8QG3+U176+#1/7S\>M;7ARNOSYY<.B,7.Lb3=.3?D?LUg)7&)AVcK70
Q8(&&5RZ?^XZX,Y(ULK]9_E9ffZ2@:B-b96164#B^Z,23I(YU?b#3O3c#NgXUB@]
<HD(\T-0Ub:8H+A<.O92fe>F]ZZ\aVODCYdeTOR=^RW/;RG.>LDTK<Yg^V@FbG4\
).SS&/GUb+#9Ge88-afSM046R9eA(?+31:]YWU3e#ZA?UL<P]9W5)8U9?(b-+;5a
f.CS<MedQ7R2Pc:+N_2c6D>:eB;FH4K\PN<<9].6/8Ag^HD@Jfg.;/+C)5.38SO;
N+)LQW[Bf>?8gcX@;7GTK6#b_dX&/J^=(AS)Kf0<P\?-JZ:QVI^5RHdJGZN4A2=R
D#KE@IIAfNYLd\,_J7LUf:N@^++(D0.&5.YCaO&c6YY+X_)_:=N#^ZD(T<(5C@U7
<OH\:d;Hb3@e+HG@GOC9A7V;Ze9[.MJ^-IU4G#\AY)2YbT^+dXR[B=,U)?g(]P(e
NR0HI=G7>A\[-##^5fRR=LCG\SaOgN_U;_M\K0ZE7DJWN-@3KR#]f-).]-Y&@ZEF
XG)E9)Y(\O&=MY8@DZ^0OF8&VJ[NIF)F0Ob7BK=/Fc<Db>V@,)9PWDHgYZ@93L07
66KP2E2@bf2V#8\fgZfKRZccA?]34+(#<S+)F26C.#1RHG.Tg4@EF9F>CcE]K(VI
=?THBeLD5TFF1b?;fd]G&Se8f>-;G;]_X/SW74#S/&gD#+^>2V19&Q=71VSd[CK]
&(]eaCO8;#SYUREN]+PBfT0>8SHF;,M+-X6I:SM=K0X4YJ<\d=F7+:=3P?ZdC[8K
3LF?12EcK[QGOFH]-0E-<SE/UF7//-AScC>F?U<.1V]))1]S,))e-W9=NfV.PXSB
@=Hc\:&;/-6a@]\e,C)&W4d,NEU^c-Jg+LVbPXR8<(AE/HXIVNQPF)Z,3XU=Y+9L
VB7G?(O&J-=ZET:G[=LcYcH+8-J/D[.EHN77ZE9;@\JNMZ/ISad.\+4K?;7KO).^
5cgac)IB0@:FFUAU88Q^]O>2ggeFNbKAMS;dXLgVRCSN2=./J[M5_-371]5Pc,O.
@01#/YA8==HC/Q(8\gbEE2M;<\[B\2+_IB_JU7M:IBEZH+(ae8FgDG62ZE)_XAUR
WDU7O2F=f;Q4CIH.PX(B,@U5(G_]@B6Y<5NW=+[.X\)C_V:X,+Nd0YLTNea)W#E_
+a1+A-2K>\ZFf6IX9,,9Q]7YWEK2C5EfWW]K&5ZJCG&51ECGU&]:a2@C>VM?I//M
LU_3A/:b7IZY@J+KHS37L:EVYG=K-&]X6LT^-3NE[U7HO>#3202XE[6HEM,QTeW8
RA0>XZIFUG\0,[dg=6PBHJ:/5<<8M?aER+RS7dNeg,@/.TV\R/09CI-K):NaA,E=
JPPI#0LfYHLa2Z/#J:[dB60QGL07@DK^;U^2QI^_5K6(9;0cV>^(+3L[3cX6afJe
9]FLXCdL8590Rf&MCO6:gTZ_2(8_.LDbE-6Q4_-OW?VL5<[81H.=(B)ZBbANR74L
GZPH0bUGbJ(CCBP7g9;/QHKB;QQ1O<dQcZ/G3Q;-?=>(_(?[KTB]>Yb1<0[d\55_
fN;EF4^9_@?ZE5dB^_F<GVA\/FM]:OMLDS@EeMB3?YERV<0gYK5WW)=&:-6E[43W
aQfEZQ^R)R.]?Cc-b[BN;],Sg&dDRVGDF8W5gLe9CPC.OAN6,-O\WZZWWUW.;PR^
O0,8,4GU1MFM]6OVRV(4B^Xf9C9c&NR?2][NKX-)9689F^6<EQJ>K3.JZcSd[SNT
R&I:JJbV4\_bBIQG9DEbU9OD>6,(_O7USSESC[VA,adWM?:\3eD4KF+><E9>8KCR
).2WY#e4BbD4:e>.&0bAQ_,<_2=X[@WC]_ZcMLK^FSf#FV-@EB>:I@@:bcN?2<T4
:?NI.1?#aGY(7E,4TREC0.9N1:(G(VX7,<L4\^L+T[&1@7/[J+cQ7]_.=SO<bI/#
-4RY^6E#?J/9:Q1eFK<=Z&V#Q76dBS0S)787K.?_Nc4\@Q>Cd9KI#R.:LDHG/WB+
A^@SQ,4=LA60B:OC^(MFD/O=Q5V?Q?75TLd3:3SHe;g@aG(Tg?W988AOfUPE;8>G
_LJM::Ida_@OSYaWAA\SZ2:XA?>b(-be)Y92(/gf(]e5/EJ,/]8c?dA&,H(c);cN
b283ROM?f:&JU^[.XE00J<JWIK^-,8X1+OZQN2T6()NR7KX^58P8AGU0<?aV058a
cA750MecAdT4/b?L#00,9<U;McVED[D/_=Gd[@F__(9[(VHCL_3:2bW=Kf7PEIQ]
-gKIMY8;);gd//,1@SS_bL(&;WX(F88<.BD)(B,RQGDXY;OFe[><&a<DRf;E6(32
O+-7<LHU;WUe+S=RPJKAV,N(0RE\aJ&G+PZ5.KI2J92_)BVQUTSJ6(W@56M(Z1_>
eg&8KV3[K;M(8VBc)9&cS?9K9,EO5[WMO-a7,=_&1#a6J.#F0V\\43R&Bb.;4SK\
=fK<aP?I=50<#JP?+6aeD#-f#4,,92.WPBd);^\+R@3cCRT(PO,#8.-E403g4?eN
f8RJWYY/bS0T16C=cS7_5c_MNN<K25Rfb[0Y6E1b\MC/HIJ)HbMY9M.\#OGHV(]R
TRR^7]#<S(cZX@4\4[^L;Uc9<S2RZ3g0c20]<X=Ca>LH,23WX-;65Mf4)#4F-HE]
R1KFVZ@2cJ(WW9aQ3C2AVU1+@S.Rb&+\?E920]X\bHHPbE,QC#^S-b/NbDLbM-KT
^59NS=?(HGNR)QQ>X]U/^3+CI_M:ZH5(]cXfU)T)UYKgD)b3Q(8d(Z:9E.2<]fa5
eLV[g[#D17WVceFS>>Paa,>O0I+M)2@#PDO6(,>O?8_JA@0=,QDY2&A7VN&&N8O7
EZI>7QCd-BTCFB66>aQX]549d?C<cfL7OS0K[.UI2DIF#-CbO;g([2G:=]eTV]<?
3dB&d(W;a^VZM..FYd)3eKGdCaRJB+7R2RgJKgIKaY0O+K#^JS[@)8bQ__=K5PDV
6YJ\&Rf\P[VfdT[f&GP[:FO-CC,eVfBP3Dc2_=5E(EE]/F<9\;^aO+^=5&S]b?LR
-f[A4,B,P&/+2eZ9Ae[\HRUH).gg#fXJ6RUgXOANCg/Q?MXIaHC[[f#5Se?4:(_U
<&)M^=-=N3W?XIFJ=^.ed:5.&MPRNZ?8E43dQ;IS&<V?-:H)#b0f1QR&R##+VOM]
VW-FLK9<(c5HH_PU79V.@I_;6#XD?c5]GJP=DVU^<_@a@P6A?93Y5H57a&WWGX-M
OT5BY.64D.7cR/8YBb>&IL)5)GS>,JU7;\&WO3NDdLe;(.LBTdA=+-W<@@&79:6E
fTIMK@7:B-Mb<Db;.&g\5a[.2&.;YZ>])>0gG2KEX7TLU5^(U#K&35?SH,:-RVCT
b/b]6/E[137@(f.<S:JJ4/W=ZC.Z)fJ3:DF;;@E0AVS3-VV#W:&Kb/G1/,_+2:Re
K).J5([aaQVW,TR\WIaN@QFUU)5;ReZ/)gd5V(e/C,8@8YT=EO;U(W3[BJPLNRF.
PfcI.ab.6#ZL)038[:UR<IG_O6FO;(;R()7X4UESEbC98eZ)Q#Xf#b84/2-gA47\
a8W9b:3D/YWc]H3^>QNJ1a;V@N8UTg+)e6<:)g-<(\>fZ..B\e-.,A=QX[1Q;(C4
OIb6/]&EdLgZe/P9feL2E5P_GOWd=fE)9>]5RG+4d\RDK)#)/>V_;ObOIW5J?a)W
JXGL7N6W./FV-T=M7bbbQ3,,cKKTHLEC^dZ1g#bDeL.Ac:@@Y#Ne#A5K;,VFb]#I
F^[4C@@FKIE0Ta[J)/B\KU<?FMW)^=\2Gbedbf.]H8XYA29]#?U\5RCC3FE#:W#R
L.D@Na&,DMS;<ZBOZ(b)5-O@NK_+C[/eeQRXH?<;WA9MK_>5R:<Z5B<DSQU7;;];
^D:<-05VVB)S&(8G.a4+[8_U?.@9[gZN9d&Z4I:,PHL[NKI7Sf6B0:?9)[5M7dIU
(cK-E>R[@A(;S#LPX5;+3>3K8:>Eg7:4#=_3BKH[X=2EG94JIY(7PEG.2QWc.[4Q
#-\F;bGI2N9-2G:@/,N^<ZT<#+-68af;QMT,F&8.30/S[I223N5D.8&c<c_DIL4T
F(gGS4\:F)e8-KP..M#E#1a1aW]:X/6@UWa>0(=8JQ7^5YQ]a0KfQGSV(#;PTbD#
N\LR\;.O2<g9<TQ=(Oa2SAMaD,)d]Lbe)?R;MQIFa^(JWM/IX+]\7egBBL[>F/[G
?PE_)PEScb:1]TDTA1(C75P_/5P&YK]URBfC2We4A@8CDWMSX&78=Q9-\THdT3K9
+8@]2c3[NL8+,D-HRMGcc0\T]G>)-EXe;LR-?a3=KH>[S&UUB&DR\=S8DH<I[#5F
QeQZ9)][D5T,W,4TBNKcI7<M0@0;B:^\2KN-9KY_bVVT]6&_U.JeEA+(,AcUaDQ^
QY7Y^T-@03CA&MVDCDP=?Zge>B[D60I+/eEe1.VL:LW_N0D&=>?U+3(;2e;2b4SA
7:1d+3;/E1CCY<0:;?XBU^M8(V?WZ<Nc\F?fO1CSS.HXdA;[gVC@8X.)NDMC=IHT
)X_MN-(R/#I6:(6Yc?g0b\OPK6SR@CM[)A7YF)6IbE-1cQJ&:)//0XKW0gHLI5TP
MWP?]Ic&c6(>T,4NMT+XTOc=.VT3<VB&LZ:,.,]O7JL:9)R&)..4=G@K8=-J4_:-
bbMHX#;[)a9@cPP0_-KP772[b)&4eI2QKPM:]Yfd57K6eYaQD:TRJ^&B7=<LX#T0
F+/?I2T1NgBdd=]TCA&-D^8L>FL3>UG>bGR-2;a_Z@_NZ/?[3T3g-(R.>0X<G5W;
B+=IbJ-_g:)8W/-7OD@S0/V_KX[GcEND.[K+W/4[g+P(M_C>bB5@>;Z<^9SKFP=)
A-T?cVZB9c5^/YIBXP;b3IMgaP_PTZ,>GX#M(/DPCcA6E>E<;X_>PZDe@V_SfL<&
dWV^Qg:A69dK9EH^R#\eG\5b53;#CQ)&a>4B]A78;^eQa-BV5X1_M=,:JJ8D+-RH
O?(9G:U)W)S/d<S=UV_a-PSXXUHB6LV3g9SYG0EdFUI:5YKZ\P3>WLCO,&]\GP:-
.&>dc)F\5Afe3O=6CabKWHVa.(9,fHfIK,6+]I,H7C&MRU\=VWQO=(H11Sc&69;>
U]::FVW\^OP/3/US9[&)QY4XH<1,SgI?7V3gE>=B:cMPMX1f5JLXR(X0)8T#Y[f1
E4BN4,BVD],>21@HI)33-CcO3HaPd+Q(J,SY0+DaV4>b(KFZc4L=f=N3c&-=#\[+
6b#Gg^B5PBZ<MDK?++):SIe3BO<IdZV(CB,\0SIFB+Hf7.(SZ>9B<2cXXbVM+&8)
Q0;@a1bNbF9.Tf5X0gVX\gRf4g(<R@]EX3I)8d-Y<WO,/C.7[:O7OTHC@f2d/fZ?
JbD-3Pe3&]C?I1Q<)8MSWI(T[>/8B/BUH0g5FTYRY#4YJ.(C1XRaU.@+MR]\P0E;
gW]EIb(K\9DBb2\\4@fb^0394/bZ668UT<?OH5/+_)GdTc]\U=SGcBJcVa>=()&c
;7cI,)(/JaTJ\-^_B<+d4YO6_PQfM2J].)+QW\)E1A::PX\.QX/-=D2@:(YCN-\>
VO1N52,Yd@MZVcd+##[AJ\#/]RYO11:;d\_Vda@T@(\_=bQHKHQ^2JBA<DDbUHN^
_f>?JR?C?Q9+)5;.P.,I?8JD6+3c;F(S3S\BMZ/aC8JF^&gL8QZGH(g@Kb:\DOUf
)IedYEXOZDPJ-G?DA\[3aaCcQ4839EUPg2;J3^K;VQO-EC,b<B/Lg,-I,BHHfd&)
XB<]Rf5bD=5Vd2G3gR#N>[4Xe82Y6E<?RbL=]K+]]2HW5MO1+)+I2YP8/&RY6;9Z
e#SPa^M>1?=DP^;]La-d4C)W8bXfOW4F=0@O,A]_YBB,2]<P?ME:=5eD7LKcYYP(
:VZ65>OLL<OZ(7)]?/\f>0&.4)@K6G[R>S@HMSP([J2WH5V&24;^I6A+I<W]#fL+
cdN5PFe#ZO7Q7fZ23L8c\];NcUKD4YFB&@U-.ZMC^V,,HAZI@XPg#0R4FNFFO.FH
aP/6RTW=1FG4B_G\+-U<1=;WXLYR/Q:TI?_:fQ60)5GKW#f=M/e4(5_(F^+IIVI:
+#E1>fI3b\:WJGKT#_TBZM[d31B[J67U=]?I[&P3I\,N_ZU9c]H-D;?a6(eH0(Y4
Z0NZ&VM@g_TUb33-DT@L]QB7>dYNQ6K-\6U-a,52-N;1?NYC#[JK/[16EO10I0I@
CL897b[_,JVY)Z9C,Vb2;fO:NB&[A[00^BcBeHLN\d:]gC2/@-S@;c#E5T:+GL?O
=6>2-/J9(5C:,>M&IgY(?XXOTOQN0AOKE:;;8c_eM-&TQ)2>31#8CHHA7OW]7dO@
.MK^[\5df76I6H6GJ/]FFN&,K#HRWL3IZ;B121]5_=9X;G#89BOX(@,:A\_:@[3Y
4g]JKgNM2Xf-W>6g1AU(WDaNd-CFBPYK_;3.I]Ya1^RP-cHSNW<cAB8K/7K3S=X9
9eT1D>/VX]H_K<aXXM_a5B01bQ(SN;d.Kf)7^ICa3]7c\FZL3S<EXVEG<1T0?fCP
Age^3=eVaBIROIUEa/[I)NNY/d6,<f;KfZQ.?]HS5Q2J]6D?XggbSI(3:B@_b]aG
9=]?#bWD^7&2QN,_Z5K7::d=C1:aHgc_.A-:^cZIX(b98)5E#C(W4QKDKRPFL1^I
Ha?YUTd/ETbH_U;)Q7cefV/BMbUb1>?a:0)QU.[[?#Iabf):/gI_:YT#dEMGT.3M
-?I6+T1?d4=;E^5.X<XP,^)81\)0Y#R=B\3@HL[0))2@U42ag\K#C.(&_I1F)Y_8
@X#DIa?+JT>0^.JdS^Z2DY)#fLR#YdN3U]SGRMDd32]S:UCL7R-4bQL.+JKQ46.[
EP-)[Q(JKZgCe(^O?RcKD#(6(.X_I/(YMCc)Eg0?Z=_:=K#\I/DR]GF_\LUQ8bL1
b_a(G.[GFSWVO98#(IU@EF#0adB\0N=U4c0Lgf8T_b(B.F?],,ST<Y-WGb(&_\#U
YYPdbA+3NB72/P,Q)R-XJM]6SLLV9;7YDDT#=b<)bcQ@1gD=V437WQE&]/PK_)5_
;eM8O^eL_J&]4UCVD,M>^+<3Kgb72fQO.F1JTTG?WHYL-K3Yf9S#(VBe/2<R>,aA
XO;&gUHO\C@d+[JF_9>EQ30F9Eaca;?Y/HA&;C.</N<VUQS^V/f?L:VR5C4.W[5a
>g+b>80>Be;-CYYP+\\[Y\5GAIR8HI(#ZI#[L=F@[3YFCQS=[SB:3=Ge\^X:)-V4
J.HOYM,SYDOTI/^)Z-OC.3.e&_Q9gN##,CKg?dG+Wc.0X@b@FJ[Z]GLe=+-W=&XR
W[V3--M&>^A2]MU2g411S3Hg9AGdA6SF)[4F6JZ8bLFD=QFHLKBdO2bVDYZd?I5P
.#1DYd9\>bW_@6-W96Q7TaZ_[PX,\4Z;WN#\8bgC.LN?^;T=KX.DI]]./f4\aJ(2
ccMG5NR4aB?9?(g2UWaPbbMYb\B^QRCV<F5]Y>+ZZ05_d>C]Kc6/N\5Q/NK_8J)a
ZQY-,QK7QN2bJ?7><1S92bZ2L183UJS[Z>&V7):d]b?</_26=Ve1X+,@-2a5_[b2
K_aPfg>LNNMI:Z8&1DeS&YG/@)K(IMHF=N@KZ3dU?LIOI^)-c.PMU(>G-+bd5_RS
/K&DcX?5TG)[Z,b__OI(c^TSHE&PJ+SW\=>XUCU1FW7MU=NNCDQM1V#<b0?>G;>9
V98P;W#45)>?GLOQdZI)FU(WbN7.b2[7?5MNWXOSCOPQN0&W[S/gI?EJbWX5@6#1
(D.EHSQM[&89L4RK&,H4K\)E6@\CP3X@IEXYNa?(EKK,S.GJGd;MJQOBT^H4WFH/
d2RO415M-<]DBPA:S#-^:FXGJ55ELR:(AB-AgbO2edVYX8Yb+4,(?,(OX&7GNb[<
)If6#9bdf+4RTMOL)JIa+J73[HN0U5cIPT^.O)/+d_F<+9RFV/9+f_197&:?T2N#
_?0+bFG_MZQ]]H7Ue=Cf?6WF.T6U5YM\0BF1C:-#@0fY)f80JKLYgV6f@LM?VV::
60;EI1JcI>b\+R&G8=^e22SVN1Y7(&NbWgSaESb^F,Cg]SA8XEMfU5AWR5ID4CA.
fTA@L74SbC.?UP()_BGKgW/D@:Y?\N[gY<YbV:D98-(N\[\38Q_-_bCFY3QN#-Ae
&\GOJ(=R_6SL^ZD_cTc5Y&_b)3DRJDF4SX1&0g8(IDTD_V3Y(V72fA,cUVYY;6g,
#B,8E6-L)UC9ZYIA]Sa)FXS:<;O(=V:D<-U;Bg:#&X<?8O,#DFf-MaODP:LFVbV;
O/WId^#cR9,8eW_<X;P:F7<(H@4b3LXTZSMO@OIgOLN.(=SW;HbD/TWVb:UO1ZB)
A?JE^#L.3FU+V\VG5F=K1J9_K5TAH/1&@=349;]:4B@Z&,SW\c_P,eLOHH6EK@c_
^@?<^P3bEC&]94OCX2+5,c(FKV\]eS2BD#@DE:gfW0XT#[DUVP]@-XA@HddXK4/I
aOODZP\97+=WV)9]dE#AM>C+gS[\Ib\5c-Y/L#WJ6]<)b;BOLaLgM6UY@Z/@d^#H
2@5fZU@5HT..e8EI5:J5P3&56OGC&8-0B\19]cRDITeG(;#g?&6M1<>K2dbC>D[g
YQL,)eX:AJ34&=eY7+(4DZTcBB>1)9)H;QFM[0\&^&ccgN:GD.c73[M#Pg-E(HBQ
UU[F9S+OZc<LPd592bYg1VF9AJ/9DQ=,U9343WSBMOBLS^[IGZJXN4b,eX1I2BE;
RY7D7aARc9WHN+8c?DARD=?6GL/PKOP\#F43@))-3,Fe>S5P_F(dBDXH2g\U-BJ]
KB<ca]:ZQ-(f^@N6LD3.,TLJ1(2,)T5MD;<[Ag>Bb?]D_PR1NBUTL;P^B;YbMW2H
AE;cWR72N.I&06]OadVFbZ8aS3?0(B:1I/DU1Y>C:Bg_K0CaLRV=/J42?CeX7e=M
,>db5U)cWW_YQX?LCfM-Ha>R<:/#H8(cZ<(<Nbe>6((Z#_.EVH4b+Oa+CJ>D@aAY
8>SZC:gQK+>XHd1+b=]5d#(@Pf,fZ]]5CcdQg1@B@I95L.[/]YO>Pd?Cf1b@<U5Z
Z5.[A^OEI4AL1\HZD/WI<R)^F-)UT?YdVEHT\EfDI>QZK?JRG;SJ9Xf@)Lc5K=Lc
RL:2NNF9(&XaVUM\F?JT1Re9I8bQ,ca>@Q6>8af3(,PZKR\7U?Eb+[?8L8ZBA[HX
g>KKaH6QG8#H8IPWGHC)fbd?Sd[.998TFP5RNW&,M)XCK;WC3X6U_JR7\^&TK,EM
Z5PX0)-#LfE)P^\2/4>6X[Ed-R3AF\K:LB-O(f=Ze.541N_Yd[O2MYfY4ZQ<>FL6
3c<ge(4^Q3KF95fgG[>d?GgE2e)]>R#TR:f@@/0Z4:HKG?_Y4,9IMP8AcBYeP^c=
+MJYB#0d&LCHJ,=ZYZ9#J2MB+7V05IRQgaVQE6GI&D8JGUS0A6S&8Qe+9P-gb;2#
<K9Y(bI7EIKcE:]Rd;EJ&d3&D]0d,Tf_\F\7M[2RHT^0U[fA<_eeb1I.3YbL1bJe
WSMRd#9M0;/,=IF)TBUL(9b67)g8^.T4LcN(f_(A<gbRW&O>>-Xg7,=M6Fd^8Kf7
((e0&/Pf7;HZ;#HYB+C(STI(B.5#b2I/E3KP(NeVf9+FV?X7H93AJB3@+AL<E^?C
+0[4+?.8@P)e/>^d9:.)b?6+OH?)(g&@^6eWB8GU[D5K_N5WKU@P8_FNF:C1I?:[
,>20:#X9Zg^IS&-JMA:CNaU+g-(6\EJ>e+VC)Ia;Z&RFGMCbK2B(3+\_7SNG<C&<
dE13V?TS1WG\T);W+QD^79a[]@#V^B\6P->13HH?4R^G?NNH;K(F)I<K29=>4,&_
)Ya,eZM/eD,:>F=^UG^BE]Y;2:^Y+&)eO?]]O-bW>F[Y2g5(CWbMHC\8<@K_SKL#
3/dZFS/MZ?JKc)^Odcb;a2?D)D>(43,\5g))b(QL+<GAe&@b[^R4EfHYHcZeF[O2
FaA0/5>,aK/)0]a4.V4A=S-0<@5KN-KLFFK;?R<[+aVO2:#HP&;25Mf=cRBK8Ad-
L[e0\^3,,)\EBSb9AF\R=f<B02?&aA59>B2Ec:0^c<T(2);a4XfGENg_ce1AA?;d
fY.3DO16R@VM+=<?@4/YfPb0BK9YPY_C44IPS9C:X.C;D32EO#JY3XJ1VW;N3W8(
/6.N6C@F_VT>;Sa.-2Q)MEIA6a@A2=Y<bP;2]0D@GPc;(2LbE.dK1X0P40KD,2/e
E&bJ@8)GI;3_.JU+=4C-CUG.YU3a6[N9+P<U&#-Nc;,(=Y.Sg2Z<[=@05.0MZ2Rb
fSf<7g-IaP((BX0\<T?CC=O^P0W)UHRP@N9<MOQ)&0H42Y1Pb#X@/4e2B_^)^:[+
465^P5FU<Jc3a+f)0G:(cBK(U)cYUe&9@4_=PI\;,,_2&E9cZQJG=#3&.E8ERe-g
W9(NPI?NG,A>S8dd2@3e;?_9N:@[[:@UeR.2X@-a\U9_A#OF:_dHNFJ2;5U=I9\b
7SUe@[^c^+)/ZB)a7cMG@K];H6L_QTN]E@<)8?PK>[,]=5N&cX/M)+1@c,Q65.+g
/>3N4F.?\XCQ]KQ^VFa^W#IaR&@]_JSJF@f^HR^EBAO/@]R];CKJIaW6RT(Q@USS
Ga)RK[L#&_.SeQBA7VO\<#dcN332f]X(gW#cG_#(:GcS8bGBe3HGddfNg)FN/9>C
e.O&?TJ]XMYI(S=T\V-Z5<3@].\/GH<g.72\U4Ze8+Ac>#1J-?V,FW<g<6L#eZEB
NTfM17Xd5Y7fZE;#cC]2O:E[?9[U>a).-)d__347<>-N9.B>=Q/8fc1@O81RUe1d
Q:UP&6dJY7Cef8>0;<-UU(_(@WHJ(N51aC8\:c=&\0@6Z#T5#0eGI6HVc2F8gJWJ
>C-:W2K)4;2)T063F60-8MY;\1=<B3,cbKL.6I]E3Ucg1;b9-FMJ],D(B/S7E]]2
^e<\39E#)].H553Wf\5fY3R/#GDc-W,_Z@L/TPZO;AC\H^]W14&.5=8]RR:]M)]?
b7WHee0SI1;<fB[I[c2If1#V/5(^aK\(S)A+E>bc.#^8XO_AeJL=)H4H4[3_K>g^
fK?=YA4bF^)32L301Tga7Eg5dQ#HQEdDU^Q8#[d_?/4[42_8gU?-[b/=<H.[N9K;
M@[SG1M6&4+<4g24XJLX6;fF;7B_b--KQY4_#08U-:f(BBRF(8&ME\f[II#Z@55X
OH?:S4/-@eNVbgbGc5_L8?P5d@:W/CG0<>;#H&ZB<N;e3;#Qc)5gH9[=Xb_0I8U/
@E>YNZ1?+UWMXRYX:M6a2H/D?@O.@^IR+&^0P-DU=95<JV(^fGPE#,YI.7>C-5Ld
LBNGUH-L4dW=TBVZJ4--P9^6-VZ.45=<MRH-NN]/I,6B>(feJ-QM5&c,AFa3#&@2
]8>b1bf:<=1I\JC2b^FJ+QcF]Ta/:K0V6ff2JHD+E##CT2a0QOO&9>K=R/Sd^0?>
Y=DbHg=:8HK9D==)H7Tf3a)WYe&?_R)+]d3)3La5c:L#RPg[]+F2K66R^SdgFCX.
.3UMb_N.8.Sd&_PT7<5LMX>JB2#=(QOFP=6fU6Qa6OKX>=PK>6ARU0BAIBdgH0Bf
6)VdK&W^[FRGSFbS8gIKB;C5BI8&C\&.EHd&BST(IB7a65]IUK^F[6:TC;=d58-@
ZP/aD.LW6_f1WZ>1GY[GQ9GaD+:@;,M4&OG:6Q+NCgYdIS6)6WY&JQF+2(,Ub1JJ
&:T1fV45:CWAWLE>a0T@Y\53OQW<D=2(5<QGa_OIZ]Uc^>_GWFa<#bV]/(U7\OP\
P/cab52GHCfBQ4+LJSLgb3ZL#CTS111WcPD7[&\QV4I<Cfga#<@.c8MaT)V)FZ#V
)=T1EaGR?W(UDS_YBXRE:&,Dga@>IK6\?g]/MMDe-9216I&c)[fa2V?.3M:-#b9=
N)WKW6B9#0P^[F2A]#S/WS2C6U0+5X8^Dc-0G^V6GEU0S)aE5_T?&0eRR0C<:d.Z
Z4X_(4D=X54XZX+X1,0gc857+RK?fT3Uc&4c.&]XdgaJ=.I]Yd+d7>1bX5\C#^a5
Wb_7@/Yag[]S;2DQT@#HYB;@)ROQ+,Zd/:@4&>#9=ST=\=,X^GJ36Z:?T\7?P.1f
gS8/<17BIS;dZ8ZC:?HH3K&IA[GM7Q@AA/PU77NZRTc,W.ZVA8e,L.SXYDZHZ<Mf
XJ58GbI)\75S)OL,)9=\L=_DGGUe,I\LWYV7,1QFW3GGRQ0:58B3[_I\.(V-3G4:
c(<?aX9J55UJ7VM.()5]/9O176a7\f]g#7?;GZC))\<e=?BL)7B#<4BCNJ/6ZXQ4
(DfXQH3gJF#4V2MKCJ-E.01,c2<A[?@Y#@#<@.#<;O&-4XA7^MNV^61^G=ZV,E;<
U>&0dZV\^1dAYR:(c1..PZ;XQ3=;8^1d;H0BT>ZUS?W_,J6(,JNUEI0O_fHIY?H(
R9eQT>_cK\I+=<F-MF#XaY+C[U+Tc02f.^K6=<39SFVSLFSM[Mb5(_:N2D<#9J0T
WCbI<KLAbR^,?V,9W(<a.bK,\=6KAP:2gOTV@\6;JcfS;FHeEZ&EX\<Kf,N>I]A>
eeNQP_7bULL2e8gS1:gK;<O0F6-Ede@8X0HA)M>V):MUgDS<YTRS[d::S2BBGV&Y
UKJ([W_5GFNe_:#NHgUZ8W40fLL2PF[BBgV-?.C8;2SC>0L,U\b6/:)7dN22Y.-)
8/B8LdLPK[1OgQ,8)4Y/#MfH[-1ALaA<cAf#+bZbO[AL0Y;3aF]]P)-@)?fd?U>/
Q[N:++EO_)([H3V1XZ1;2C](7)],2C6fOTCJ&gFAQ]ca^G9aPGK8\Edc3L9+Gg[:
HQHS&97DTBQ__T->7/c4bCX80@T5KQ/X(0P]&/6G&c46OL9Z8bK-;a7,M\+AQG?L
_Qe0DfFF(/A?I17PF/eO5#9CP;fPMZ=5+02C0AC/9HWb:c=6+^R]0gYaT#69W.-V
A<@gA>^c^:G1AaWQCB_^U&1<ad&59K2TIE,E(PRAd(-9gGTFXQ)?0\ZECeQE:T:X
MJMM?2<^&\/e0,-OfV;KUE<_If6Q6Ua0CUY\XJ-.KCG&YSEQGE80YJ9e3-^8<YY4
O#dUK2[8B)(IN))VB\->fD-?)+?75HB524c@UW-1F/7b+/+/M??6REO&G&3[eAN.
TIM_<+ZFL+0.)];IgVc5-G4&C=UM&UB4152E5[Nc>(II3bJ-^KS3WKY?=W6U@X?G
=IZ[PYc_LQ]?,VHC:ORO==6925YSY&gK@2aeHUOO/V&[#.b6XVG^UTfG@+9SE=46
g(908C]VaJF92_(QUYX>5g,0#=LJL>H6;ZTg84L=ETARI/;dbALUb\()AG86?9J<
GZXcGJH5=Y6A]X/gGS9)M,KQcPM@<YTHSa=VDLTScS8bP2RTFZg\E7^W=^3W</E?
d;RNHb4KCP3MPSNMg2/&)R[^IX-/90YP4KM7aZQB^^F6I0]GX01SK1O:3PO1?T5E
F4>92(Q(3af3-PP&W,c#R#(8FVKf=/^)95<PEB=TM\RDe^A([.O6bU1]d4Q4b3&T
H@8cC)?03T_^4^8:RaL.]E62bOIP8O=3+.V/Y_I?PP#IU.VU=EHA4D?b#aU@=;V4
1JPQdJJ+]YgOQ@de5f7.2+,>ERF/]0g(G]_E-NQ2=ee273@;+;&/4C1SU@f<VOO=
HQ06XO51X>,N5:WWEWe;#]a&03W[6P857f5SY^cC3If(S&20-TR8;8g6aD88OL.;
43ACFZTM<.9HbGLJ:6+IG4d>X.9ICI4]WIb97VcUf^FVW<H#D2^MS2IgWNU4AK;P
)X(eXT:VCMZ5H+/9Y&Ng(@.Fb(2R[]>+5IB5ca8XJ2b+FI]PU;_K-ae[Z<I2CQ-F
eXBCKWU[J^TUMbba/CK-/OG^0>I_I&MDQ<Y)>V[\MCW7d@/U\#&;^)U_(&I<3@gb
_GNOM[-VT_0eQLKK[A-22e<d6bL94=3B3/190_W5+;(;#S]JBU1JJ[[),?QHT_]f
14]Se_\\N&/=6+O@?Z-DBb[+)&&:?Ze6KUb[Vb.99.N4]X+gfaNDZRGQMFg\CI2,
0d>8@DLb#NTJ_H#OO5\B)1FSC25#9,IfZEE1]B?-e:[g3Y]-LN-LD5UTEJ]3EBfY
O[)>[9Mgc.Pf)DEWYe+;/3Y8_DN13NXS1D0KUTec0:VK^J^9L:,e\714?Jg?XXOZ
\V)a^Z<f4#,:.g\<>e4>0>XV@D-Z8O@3K\?,ID#6U1@L^@=]9YVFNa)#_P=PA^;X
J(cgbTI6/#:.AF/Q-HF66#c+fN:WBI/B8&f3X]\\BDYI>fb)5gQC.CC6P57,#B15
3<a<,dI4+3P7(,BS3FPc<VJ](&S4-)/K4^)SU14EH(Y2Q(E949g6T9:8&ce-OeU)
^JOO6f,LP4OQ?\9P<#K\]4e\9:cYUYCUOH(<R&RG2L;UL)]M9I#8WLKZWVWKMa5b
@Q/7EdL,SJOaT8;#E>>J90VGaX.-.251DLNGOX4WN)Q-O9[Vd5>b4^FZ-c#ceI@1
?W^c6^I<IcV[;#X0W,M+7d440d-TQf;:HeX+(O@0;9<g49><VFO8=.fCCg]24OFf
]J;8VZfD-[>C>ZWH0=MZfXRP4Q]V4e2IU?DLX2fg1Y-VSPA>RJcb&eS99:+a2dI:
L7SD@4W:A[7WEYF(cXV\5]KK7=8/I:KE.;UTS.a@U&g>01(9UR1+3J;MPX1BT4>a
&GH@0J&.(>.;5/[A_O.HLK9]Dg6]aO]1+c>M=Db\C..Y-0Y6CdGLFKdaW4:MR0:]
B^&#GPg7PCML?,.T22]=).2E7V0aFXU_BD3@_&I=(a:J-DeOg(O&b1Fb?23C]2TB
(I1Q/T.JfgRbZ_7FeA2>Z)S^.:LM3J\1R)?@4bK-/dEGX5WZZBOY>^a2I-H\4-Ef
;(;2P>a0?-QEdL42W;7IbI_-MD5J9aN)1.VEeU:f2bGRQQEdM1C^Pg33SZ+7Q9F7
@@?ZBO(;9#\JZV_G5BB?@OLC;(@(L].[X3Qe)6GN@#V<6BM#.^SW+,?DYMCR[_-b
5N?W6,VW=]?HT0JJ,e2JZF^2WWbSGRa=:9:WC8c#5V/H=E/V&OT<T?:8Jca4^1-U
EU0T<6)aUW).3fI;?[YB_I5Wc/cc30#+[=CeaMaEH&.4&XTc#MDE(;RM)ca+?3c?
>V;(Q]9bFZ4)LWb#N<U<.#UZd7PQ,A/QTE[\;0[O[(gMFDe2)b5Lg@4#>170C)-T
d65>.+EDYN<[Jf2BeI5M3\)S:RbT:#2W5R7I07Q.c]5V/G.I;I8NFM1aF++#)Q>F
;3S6H@V\>^[P7e<<A,\#G5ZR+XU[:f1e\e&cNNL/;D1?FLBYD3P?GNKL.^RDPDBG
PegRM&9/@-MLFY_=R6M=YL2M6@b46@>B[H\N>bK1A3>aaX:cVGJXJ-WgUW.I<=5V
2dQ0FT4QP^>f&BKd&,&.Q)f25_&[YbG0?=]T&Ib1++25JeF/0+[GS<O.P.9&CgA(
8;T<0H>J<d;?#O?]MVM;=(G;,=-/(MD7_C>5;W[\X-Fa=BQ/>ce74?f:2&W/L;LA
I@FS/>-BW,S6EB_dH557_0Ce@X(]OYP_&>F\0++=.>(^?MU27\Z+MC/QU1<\XN?3
DJ.82_^[ZRd@QgFW<,(UHDD+__AMeEG<)3_?)]a0+BF5N[(5)3C3+)Z>UVH-_e0O
5/QUaS#Q8[SH?7eY&G@/JI2E.gV2YG3D5b&bNZbML(3VfPM.G8S1T(gAAH19-1?,
(G9PJ1NKY+e\EWBbHPRgMOe_]1P;S#dRY)eQO4/JID@IDfX2A_/JNK+@)@G8Y?H>
:/>\[:.>D14Ve;94&#V^6)\2#_eSg3_OY^B^(Gf6#<)cR_>W3G0^O8VJEOaW#eX-
LVGN#]B6AG0XRFgP;(\W]J+E2DM1\)5H97]9V<dZ9<RYM95\+@&EQX=:3IWG4::J
4^4:g;L,J+(LA1Q4##ERQP]RbH5)B&#K2GYG[8e?0X[0N]<QgD2\1+1142<KR[:L
O;]Z[<M0Q=NK[HT01,T1P\Uce_83KT,P0J4-A:5aH\Q4^XL,M-:EA&5ACR->eTVI
63D+-AKEWW[[7A=IMTRUAZ:Rb7#,&9JCK?[2feH\X6TcG?LPc(R;c>P^fF-<=IBM
+9ZR/.#cOXOLI50aV)G(ZC)BVNc?.74>9G-SfA-/:JOQd?E58)@,8C@I:,Ad,H7d
+eUcH1JSEdBRSBWK(BEP(#N@6BCT\(@5#YTW9D#IL+:VU4Ra@OUYcXHU6eK[&:@=
L_P+^@^HgFC5gF;H\+4&7L>7d\<])Z-M34Y2@T9NcJG1cKDU3V0SMIe@(>-\\f:1
+YQ])MGP;dWVX1>B6MdS[/BNM:IS_;;ZUOHDOK#9SZFJ)][P#OGQXC1V<Z+HLLDf
fdQ)EQ_E7N72S#bK])807/01QH;UW&De?=cK,KC:V8R@c4FbA?f^XPXCN[:U-]+6
NJ.H_,4X1CM02ATSbF:IZ?VG:.;VQBKV\g@5O_Q5U@K7W[,a)//:@:;bZ&gYDB.L
fc?f;LFI\[M=B^DH3&.FTde0_Hd_D\YUW+Uf-PK7,^3-YP9+_FQg:^-F@R]WM>N\
c7(F#^RV8M4F&SbL[AJFg,_>1OGZ?^#IJ#cI?3[PUKGZ.2eQ;_(U(f&]\ED1M^M)
9+MJ/0WAdd]/R/Gb2O-IZ.e9c2Y&3M@G?G)aecZNXB9J#O;M^U1-Eg<\^+)e_75c
2J6Qg;e/IeD/6)P,#233Y\3#A[EEEED96OYg+^0QC?@7g-10II[]>3V-DdFN7<@c
7V8eJJ(S-:.N6H?B?\VVUO_JL&IFLB3(GO#4P6W>ZLa6faP[CS6??P9&P2H[G00<
_f=gJg;6X@3a]TG&)TPY1bI)91Nf78C6IFB=HNOC:.HgOgTfN.+8^2bbZ>Z9E;D,
SMX;25JN)8We/=3[Sa>)S4M129.8&G443R.\e(SH^KTC0/A1fPS[A8)?d>97L]:)
SGF+eRR7NV@5\LfQ0YCOQ(YPg?T&H1[7^)Pg+[YY(e/F[_O7X)Pc[:Sf(U.7+SJ=
;V/W,PeTME-g?4R;Cd&Y-)g?2=W+1IZ0/<[B8IG8L[C)\3;-9b0&-/<Oe/->AcL3
H-(O.RV)f.RgPB_YBfV4)IeRM5-;BbI]fTXW84I(K1Ke(N64TV75bE5cA(MNDA:0
L&=#H?^?Lg146V2?U6b9OVQ,Y9B6gIH)]#MZO?>SV#K::(+/U/S9=6OU3?K;_Pgb
:68+LDaeC>f=gDUOV/4_S5;_PVAc5&/daS#Q3Q#(,JF^W28dGdX,VGSC+Bg32c=e
2dYVD67TE.VR(<I+GgRO&1,:].:UI/FE<.UU+d@4X&AR(e86WaWc:_5[-WS3I^0S
gO/-<8Ad#@McH\)a:A=RB#;^Y?R\5]4,3f8:]9aGK\KA9M#dB?aD8_)GP@CX]ZT9
/0(I>QFdaPS8KIJWM[0DV]=D4Lb1CTR-c>DLS]HKV2JaLPB[(1Ng;?M:9=4#:7Tc
JL/9V.T6.FBYGFM\);Y+/:++16M-(UWS6T:(GZ,3T(./73c_85<MQ)_JN-E/VN2Q
-2c&]/UW=3DK?[7=>R390If-?KFebCD9VK7SKAd(0EUV\_5S./30>HfQ_VKc+-8O
.+[SZc0)cT3AB5DK6MFM2W4XIF\/8DG1S&QY;UE;CB83.F#0MRZF..V?_KSg;4<I
SPXY;&8TQZ8e1N4Mc@_U,2QZ?1eE;Hc2D1IW=SKY)>]dc=3]EVDK7)I(.O)cKU6c
=Z^(#E&CcINU>HWJFK\8D+AS)15&WYa0TD7?.PC0aOJ>SD\LN<_:9Yg.XEQKa:d4
9[_L+aNQ.WC7([Q)WO&.^;B6KGDLB2=3ZN2XU1LA>6dKMD=0?NMZCM8D.ZF:@Jd_
@5Qf\ZVL;[]4B;FfHcaTd0(6G(H(MD-X15_DS(825NR-LZW?[(O/K[VdC=)(2f]A
\QVMb7/aLeT);27Xd/a6(bLPJ4ISdGI5U&@<<NMFV_^9KB_W:8\6g8JSR>9C[GRJ
\b[NH07WO@59P#&?NeNdPZ<ST.J8O-X1=e</&G+Mfa\@31MO\,-FW;#&,^H(G1c8
VH_?e2L\CF_O,9IJ8Z/.eR5_;[=BB<LE+:)E?aM9VJ9fJM-ReWVE972M9=?(8/([
<Y^RZ7HabU56(=FCdc)SCKVA:Z2L[5T[6Q6Z_[-@cW7(b\HV7C81YY^DVP0gZ57S
[TEMb-f3)6:R@M9[TC]YTgfX0?B^N+[2^SUMdEWfM=02SHN?U2I09dLM_ZSY])@3
:K8gRQ45U9\1NX>cP>MW7\/(?cX(6V=dEKM-F<dRXKTg\P>#Ef3bedMT^W,=0,\V
QT+6THA1e=-KZgQd#6Dd/([e2W5E\>e/a-9?@97XQbf5@W+=L@9Q7F04,@+XXe(-
ZXQRKH9-SWC_+.7>fWD(:H?5G+AO^J]Q]@3,5YNAU2_C#@&K[fE8H_@M.6dP4Ce/
A;L+81fB?CGP+U/KM]L4&R;aZ/(8T#GJCKAfd5>;@b+bAZA?g/4-Q^92KS)?4?(P
aRf<#J_##8D&,N2I2/=WE)]2:/;<N#C&;,DbUN@:XE:d>7b^<HH_/K#GV:OWO<G;
O&f)U[<6d^6S.)/MZU,8<93]OD_NfHS1)9#8B=A.c\:MXK:ZPV,,8)7c8;7=+O22
G)?-Z)R]dTX8<1:@Z(VO-KCgc<ODBe2N&[(@cI9TDAbKX2?>Y(39U?g-#DE[TYfB
O),0dAF>M;C6WE2-.LSD9ZY>?bg:Z]POK+R9137e]_0R@F_N,aa[aXKN([U.,NFZ
N_H&_+J,EN)E^2g\N(aVV2?(ES4a8Zd38#?N>D/?N]5dB/SJdV28.>Z5K?)d2Hd+
5d8AZReYTEVa&EJ:K4HKXO]eTBU0ZaGET]](ZLI&HQD2GcVX+TK;_Cf@53ZAK&(:
7=3Dg\O]W7&++]D4@;TBZd=(</_9:OK:gY+0W^@4Mg.XJ7O?9&;H8<3=/-=67cXg
-eb3M&3<W)U&@c7R0+&D9<852I&C3>QR^1W<UbfHQ[cM5..ZLH,Bd[f[C1MedV\(
0F_+g?91d^=3?3N:g=[NFF;O,+)6EPQ3C6c-H;36Hg;<bQ33<a18N=D(S)?WW/GN
Z\_fHQ/OQ>Z\O-M9g-ebYYddH[(>c6/11/?IHTL-<^C0ag8R8[)0QG95PF+]PY_&
R#:=./fM-+dT7?];Hb=;5-K;bW>(1B^eJf=P?H.\<E)ZE80ZcPc7B2GH4C-ONCMN
3OK-5Se76.3MN8+IGP_VQM,R<RVDcaT/)()eM_Rb?/aXMJ4H?87@N35WMNd;-6#+
UQMP_KS1Ge82&/[TXHWLV67X(_c.@A+,KE1+3PY1WH]a,TYFG26+8TY2[R<bOLZI
[P5b8GJ)QBHgAfC_:5V5=_G3DOTZVIVN#a3fU&5Ig:#59g=I/dYLWF5B5WVU/5Rd
@BS<>7eSE9>I54/eI16\IPO,V0RUU9XagGRH-<FO0GG;W]TGE64M>ZV,3M-]0>Kb
0MaITK3g8Re=X#I.8V5XbMOEbg^U8G4CW;dOa7DWJYb=e[:c/&c_)HQ:)=;.-7YD
Y>1J5<RW/B&G;c8#(P1@XQ(Y4ac0G97UG]VAZ+@PZ,G20K\O+,Gc?#]H\)VBHXOL
+RK>1+Pa7c=HG@gX[bM:E,QSDc3/29:[_M,2KW/fJVXCYe[JL7E_)b9[9_HLWPZ+
Tg+_WND<^#-O0\3;e)U#QeJZSKVUZ2&RK,)7PX??VaO>5_fS1U7H1^c7ITcQMZG5
(\g=N)LQA)f6RB@AHa-),WV9W1,X-SYC=4#._^bEb2677[G<#=B_9EZf3LE.Ce4K
4I_8489fBGg\O-AH@=M#@K=]BK(HQP<RI.OL[+R-I,B[dLC<Z7?<^0;MHU&O\LT:
M9P6V2a[I-;6AN(X/=2@?31TK2:PEL3EM&0)V,RO-([EU.,2V)P#-DWDI^6<S(3S
;LeNeNN/ZdPK7aXD/XLQ-5[I/D#b++)@+^3T^AV/P\]P2DRQQ,U4R2T=RZ6-EW<)
WY-=9\NNQ>VS^J+Rf@gCdE>f#+aO)7RLN]39Y1I[GT2TRSffc35QZ7R429&Ae:]D
G4P1)0,#fD,]:SZW><I,LGR)^QZ@\<D/O<cRF^58WHM2P\93DGSZ_c0Yg.&Y/<[e
+_:cY2Lf-GD?.F_^]eEd^>FTg,0fN_L(V.;##:[eO1Ac0(:8VY[R4YL@WEJLbcO_
S80#c6R6]@K,&Ic?FX]W>d@&&,2HgQLU6N&9.(:cT8+]dW/^9XSW5^P?7bQHKOJ3
-J[JY3T9RC#_68M=<RS/ZQ]=-WSK3?2>[7BW_=-d0d1B\dAfP.96:UJf](S&C(JK
U]O:6-JC=Y92+BWMfCQGDXf-C1Ig\)9/<Q.<YU8;N._@=cX62Ob<:X>cH?X1^[:,
,XNfd5e:F0XO3L@SDg:E87L+UKK,=LH]?=]f>\C<O+V<?,VTGb7ZCU&1T1I__P2c
ANQ(?11-\Xe9P:KW@#L[A#4/e-D0DGE^XTEaCQ81V,fa8_Q6X4_>GdCHB5;#JSWB
);R6)_XV9Wa/B4>U@7<>?]O.G2E>K[+ASARgIL&b#M@Y&V;8beTK02XeM6<O;?#,
+9K;UX)_U.MfYUJbH(Md16SSVH/B=NVLcTX7#;(&W7.E#,/]/?;DS&K:3cK>=N#?
JN>-<PKge7U5?=AYGI0VM2EFZHd5<936)[@-SGa7a8]K^2O<gS@O9-T<\<9VPWZO
/N#GQVbX6Y0RgED6bH4;;1M)9(af.((cO(eT#Z<fTJ2]V\6F&N8CNeEG8C;UK&-1
FMaJdI\XFD>3fZPbM[1W9H+[ZcaGU;S\Q]BOFHgNSJUZ3&@1TH\ZCLLb2ER=?b41
28fDZ70QJ[4@\0J2L@?01)DPOf,egRO2)TU(-I]IK9WcJA),>]f:1W_>g)fe_^YE
#dY+.);b2Uf^Sd[a.a8K8C6YZdfGZdRD4H8g==TB0-Wb-Z.]D3QM]6@54UBfA(42
I]]Q025@GUS__K7P5&:-e+/G,E<0-)b0A=HIbJ7N#8Cc7RZ+AI?a6Red#=B;,W]^
?RC_(RS:Wfd\4V6+X[gMM8^BFU).)_RR\2K?UJ+?G+BWf5]?GI97&<,Q1W?LVNV5
LOGI-LF8AOF^cT&3;/VE1YPB@\=,Y]L.5VXMeS&[>?UgB/,=#77EC[,Zcd^fC/af
QS,89C1X-@c^RF[B4FX@5L52Y^A\CC3Y+F)4]6TA7><a6IS?CJK6Y@<.]6@[.W#_
5HY)B0:>gadJG.8QW\HVTgBZcIR&<7V4(VZ9Q/__)-\MLaaGDMB/:AdQ(9e9)Y?e
JX>G;LAEE+d-RYO)0CHC2F_(eD?:925^V,7J3[V1bASSg=8P&6fd.&.f,LXWEF.5
@A1a@I_M.^/L8f4VG\<=T9MFMN_d@dE=KN9<1&Bg5HWJ0>D58;eAR>;\Yg(^[Z1N
T=_4AMa2g]9]AR)1#L<WW\WU+[RgV-E[&;7->0&K=?CKB4:[#6df)3]6,GQ:E=dC
JOBR-@MZfS0fWV#cL,_PYDLc7IQ7bVcWg>Ne#7>N[8>DZ7.eF8[NUgfR[VGVgQLa
^R]8(S?dU#JNgd9PXG&T#KJ>G@gI0gE<OHNDJ2WT_a8.,?0UC4\W_)6:HeO=:Ca)
OB4g96PL9CX]S)SCCg[J;BgWa;.D4&P5)gZ#A]U?0B,^ZU+EdBQ@Q1C4),H-aaMS
LPd\#?NC5BKH@V8\.<X9;e,;1aF1JOQR)5[WMCB1^6]-,XQBcI@+B(\X61.S(5DX
O^AQ2aVPdPN+VLU1C;S/)S:F+gD&_gM<I[-;2,c<beLJ0=LaFQb/]NUb1aI#[JIU
Q0RNS;F9dH?Q9N<+e&[B.Y3;gS2#MV9PdXcP0(-^483^(C?:bZ/7YgJ).c@fUd5.
O,=7dTB9\YUM7/+LZ[S.;dKZQbA=O42g>4NOSL<VU?aR8c6P?@M30b[MKgK<aGTR
@O2^Fg9Wf_#DbK&@44dO9c0@01\d0R0;=9Cc/=?O:d8+[aO,^D4+2VCJ]PAd5/6[
]<<3.dIO#b-e=[FUV?N@[RKJ<a=_Q>0FNQc-K#]GKA:J3@)&bf=#afK:<8;c5P5V
fCUf4=Nb;OQ5PE&eMED3^aPd(2Q4RYB:R7(:M,dGM87.N.J+F6E<a3S@;[2G^B)C
>_=^,=L&Vf,UX8YNAc?1MU)8]G&F5<Y=@aN4WafVP]A-Jc:H/<aHbZ5c]C..K\?B
\HZ[]df&d4f#I/=63\UZC)P78<3-@LI(d>5:29CCfSLST[:1HT.b()6L>=RXEC].
HB1<A1X/,IV5Ha\DeZC#fQQBD\#Z[W<e.c>ITBZ5ME&5g61X&8U500Bb&#&SVQX)
W_989MHOXCE6I\J-F?NAX>gfc6He=?@U#R1+EU>1L&.N:]DY#dQ8?8B9+O=<a,N#
>]<UeOZ=2)&01GNdegY(e_,g&?e4ePEJQ[SMV#@1NXLAGEJ5#QUD2Q#(=9=e+bC,
9_.SB2FbW(55A_N3db_66WU1P1RbF6KWM1_OO+_N5S(ZZ=VV;M#Ee:<MJKM0<4NK
,O=/2>,bY3)[e-9MfZX>8H<L0Z@1Wb[g;Sfe[a-c&c\6&>:YEBV^(UMQ.CJ]>(>-
KVI(/cYTeQ5[(JMSL2Q-2fI5>5(9fY?-_5EOfUX04=ab:ZVS.0e7&2G^Y3CQ8NdK
bH<Vg4M>ZBZL>,dga;?/JY.+>[E:Q]QX,@S9(C7LGXTL1^IYUZF0_IKE8)98YZ::
T#CF7RgET^1C?([-ce]gTYcY;-1]eNGNdHg-Sc]dMRPO&bWT#cW:3+.#7=O<ST51
ILS3WP9.99?IN,K2;]MK7eZ1Y6E8g3BA/SX10]G(,=g,^2HJ/,=+X2W(bREBXMK4
a[9FK@4665CGJ9=4_M=eS@_?##1+[J<#H/K2DQ8?_1&(3X+Sb?e&@E)6?daAW^=B
AVW6#VagO.1W;FDNTI9IE7d.<F+UO,>MLc=L(RL3#E0.+IN=U=W.^<V?)@;P&gKC
=/_e_QH/P]K(WN^W?KBe/PS65;3)gIdR-<&0DdJYcf^f]AOE0B1O_)F9)]8D&TTN
ASYIL#B74W::D[07[Gb0>A?7@=1@=>;KW2a\P,[FY+Z.B>NOg5<E&SRDDQX,KQ5U
\.U(W/B;>3#fD^g>9ZO21Q]],bAB;@8Q_OX0HYEb.4.\eO3CYRPKE,;R,JA6Re<1
.@7_3Z6gcgA;7D#f-Be&2BL//a-JDS7MJJAT7IZN?eg)10J(GAWf_;O,(5./5f7(
c-1YQBc@ER_DgPfH<,,+WU6KEP/4)eId(4.(:_J,0^==C=4eR[e[(N(FLWY7KIQ.
g8/Rg2R3:X(7;Y-Z=>T_F@H/2?SA.U1R0RFHL?c/c81;1T0QIILL>_daT\=D^:J3
SbQ__>;>c]gYH(=3\<]->7;]W/8_D<]6&,.[7_EOC=V>GN?WdZY/8FB]A<+Tfc>N
Y0]-7EA:=d[:7R\I]dD1:P4dWd=FFZ)I5K2BH(]OFLGAIYH2UYG2T?IV^ZBfN./\
QX]I::Ig(,+_)PI;DO[OgR#A/AcO.g2SUb9/]3B\3RcW\D#TSgW]7I.)V:D\AYFc
#cY1F5[7U2->=ZP&M&.dF4.IgZ^f/egO55Kf&A-3P<R:@^U9,=6=J+3M-#a>g[46
]PPOITGG3\4F0LPdD^)N1N:?.\=fQ#TYIR5g1,dK&92>1W_5(ed&=\WG74@4Y@e^
JFEG&/K##@-,&8BU[O)_.@-UG?>[Nbd@-7T5I(.17ad0;=CD1<SYg-X:9.C7<#IW
JO.CI<IZaL-H(=^,V#6UUGO2RM.fS2_MKVGe)9<\5]GRd^M-G]9:T+FK+ICA(ZXe
V1.V;f=>?V-><cN2H&?)^Z.?T23g5)>>IS/8HF=T3^YbOVJJD+T)(+A^DF>9U6gT
QUZ<VB+<,M\:f8Kf?,H/FW=P_=_^M_<gKU#d<1S^Mg)D\/^aHJR-C,Q?T7I:PEa0
&,N3;IE&7.62d@/E]7R#88Y#;8JI0.LNR#,;S1(3H?.@@Q74a>;2Q9V6ba??,f1;
#9M,OQ0U=>V-+3b/K#\.WUPDL12?V(Af#=GXe(3LO-+L7FS6KM84?KLH@,ec?V-7
(aH&@ASJHO79WOPH;5:Ua[;LBg6V0GL>79\LI:c-L_KN#7@f=-E6:4Z<@FgWaOQ=
4(O-5^XG^V(JA])3)3?X)ULBS9/CUTC-,f&VSPW4/,>(8GW>\8Z\\C0.EA6V&fQ7
R87RfGHQ^aW#;S77O1>adAKVG]eL=#g06>KKGNZG9Oef#>GDAWGEZ+A7W68Kf2VR
I4-[,=:E+[G.cV^[ae+2T#g=>W-HS4HYCN(gdOV,+;ZX-O012-SOfKX<R@]MC6,(
@::\EU32H)>#J49A)4EE#R\&Jd6?DJ6a@UP([9>:-ZU:MLZR6Tf=@DL66\_,QFUg
LG(R#?>_AS87]1WCM..ZBBQ^_<&:QZ^V3\C3.OEG8+[E?20QFV3?^32#c/1?[:4?
G&WBd+YVASLK@4OfCE&B\@QS2e;>Y-2IA,#XV7+)Q3VY/=3/7NC3I(X2BM68Gd#^
b-^WPNQCY]3RX/8(-b?VM8F_@+U,1-7[+:C,;ZXB-Q#X;X7L5WAf,FK]8D(5)G^U
-)(e/^E;&-L72Uaf\LV?^f]VAU3&WL81_]N[-eLP=49UTfaAD1aTK.AFL/9MBf[<
dP/QN_,@,Qe.4ff0R?CIJ:c5_,2f+J8].\?QGKUJYO)Cb2:ZHT7HHI9ISEDaf\ZJ
BJR@ZbKe9D+V.[GXWeAZ[^P<>@a(G0FF;0f1RX;<1F&F(CG?K0YaJMPNc5Te7Z1&
d7cY3c[62)_-JHg>TXL=7e<NDNVD0g]ZI,YL;aNb(8L\O9IKR[Hf&H/d30V;1&&3
#,L^85-WS?)/,(LR<1G;4G#PL:Sd^3TGD&?dVA=(YQb0K5FTcFdF1+9,ca76PD.)
7PXI1?0TA18bS-N1P=,?6KGg>F>,(0W3=:WA^3<A82CUNO2TA)F;V:ZFDU:IY3)T
[]/W)@T;.W[4OZLU6HPe0EYeWNfS6-1OS#OZ()PTfVT8)?@g3,?1<>C4HDSW\AU/
-ZIaG5a((E<=MIIbJW)I[M3C4=J/#3@b;ad5.<&faFD>-YbUf758/^J,gF,)LgYR
T6(R._f=1b+.[\QHD,,bQ=JT[[:ERF1.<^^V#8AS9^;I)>7S/?fU(XKH78A-TC)P
\88=J.?dBEe.Sf2L:&/S\EUY[aFLJB)N)FZY?GOWW4?6O)T840:&Y:VKH=4E(:6Z
X#<LT)V1_72PYUBDDZ=[_9HbXELQNT8&[RO]PfSN/aS-EJN:06BJ^1F<Ja[919#8
Qd_]GX<,#;JO=C_T+aW>(bO[0e#]e_,g4.]4g[]#[GU^+I\NA=S>.\a83C[.]NQ;
.1>)K/NbgGKNAC3S6\WKDW7)<7#OFOE\<]C((9BHT<.:N#_X#18O<CfO/5G^G;4Z
OKaNGQMe;A4W2?5Z@M^C1#O-6,E.FH9?gHUUIJW)-&7R_=IGfJYU@&7@#>;X,gYJ
W<]D5>7Ne5NbLC3TCY(\/JeWA:7f^L.(/7J-4-OQCK2^KDI83H,7:6Vd^FWQ8C^a
]J+OeEEWG3Lg+S_P^8RK?^Nd.c^UF,Nb10?M/3SN3>&TVDgRdZ7-WQ#Z_UL4POU9
D<gDg@W]dPL+A=<LP[eEOg>N9MUZW+012H&=>Te/\5B_7L=C4WB4fY^ZZH=WS[J]
W[8.N\YVKEF-=CINQ0PFX[^0eTFe03BVc#W(-f@0L4GAdTE^3=2[ESR;S\Z\&QB7
FAX7O52OBe?]0G]d[Oe[ZR:SKVbZ@O,E=IW<?^)=8U(J5XTM7_,:F/Z/@KL/b4&a
O.28UJ[+[,W^_7]??Y7IQcE3SYK:,,L=_P6<6O@gFC/.O_@-Y,VP?c1YFQ>6/#NY
A8^GA26RXQ254SeFIa1N9/]/<S9/,.?R\-e;QdDD-)95Y)7dg4/F.PS0O7M(4_;?
A8X=IH>BLSd7-:D_:?+E)Eb]P3WT_7>4#+Q+IU8@6\>#<g/f.gcC\9g>O__48a57
/CHfM+/>:,OOaSM3YA(9;&M,VGQd-&;a+^HW[0:X\_Ca_JEOCILBMQ9SfbRI1P@B
Wa1,EIg9QePV6+d;NV\(dAMF]5_egCg<)SUY@\gAY_>:U^[/YdI]MNKaTdYaMQXE
NP;gQSfd_e1Y+Y5]/,X7N<)]6cKc<^4PEPCYf<g-+d7K89H+He-c&e>fTM<H2KN9
.^5RW^>c?<RLMBWTV1N-e+EP]2dJWLV^DQ=5=e][WS7.1CA2O&]X^9W5;JW1#X+8
1;7]<Mg+D^<7_<[8S^8SDg3PWe&1DW)E4QeO0TeM6?=gL>DBa]4HPFFg;);_#Rg^
]O)cY-I_FZ;CRN-5Hg<^SJ:dN@;@O;TJ#f+.0DJQS)UV67<Rb2_MW(e4-PS4<Z92
e^[fE#>FcBGO]g^3:-V\Q^VJKBR,e2<]BT#_:1DebW_F:CEY5gZNQ0T+ZdLO#I;W
#9HE@O3)3327]2XGRXR^\?]3fY_e:dB^3+;DR\XF>gX0=P#@^VO93:cEQN4J].7<
?G<N])M]Xf[TPD_B5B1J\S]32$
`endprotected
endmodule