`ifdef RTL
    `define CYCLE_TIME 15
`endif
`ifdef GATE
    `define CYCLE_TIME 15
`endif

module PATTERN(
    // Output signals
    clk,
	rst_n,
	in_valid,
    in_hole_num,
    in_hole_suit,
    in_pub_num,
    in_pub_suit,
    out_valid,
    out_win_rate
);

// ========================================
// Input & Output
// ========================================
output reg clk;
output reg rst_n;
output reg in_valid;
output reg [71:0] in_hole_num;
output reg [35:0] in_hole_suit;
output reg [11:0] in_pub_num;
output reg [5:0] in_pub_suit;

input out_valid;
input [62:0] out_win_rate;

// ========================================
// Parameter
// ========================================
parameter Path_in  = "../00_TESTBED/winrate_data.txt";

integer file_in;
integer pat;
integer patnum = 10;
integer len;
integer counter;
integer out_latency, total_latency;

reg [3:0] hcn [8:0][1:0];
reg [1:0] hcs [8:0][1:0];
reg [3:0] pcn [2:0];
reg [1:0] pcs [2:0];
reg [6:0] golden_win_rate[8:0];
reg [62:0] golden_out;

integer i, j;
//================================================================
// clock
//================================================================
//reg clk;
real	CYCLE = `CYCLE_TIME;
always	#(CYCLE/2.0) clk = ~clk;
initial	clk = 0;

assign golden_out = {golden_win_rate[8], golden_win_rate[7], golden_win_rate[6], golden_win_rate[5], golden_win_rate[4], golden_win_rate[3], golden_win_rate[2], golden_win_rate[1], golden_win_rate[0]};

initial begin
	file_in = $fopen(Path_in, "r");
    $fscanf(file_in, "%d", patnum);
	reset_task;
	total_latency = 0;
	repeat(4) @(negedge clk);
	for (pat = 0; pat < patnum; pat = pat + 1)begin
		input_task;
		wait_out_task;
		total_latency = total_latency + out_latency;
		check_ans_task;
		$display("PASS PATTERN NO.%4d", pat);
		repeat($urandom_range(0, 4)) @(negedge clk);
	end
	YOU_PASS_task;
end

task reset_task; begin 
    rst_n = 'b1;
    in_valid = 'b0;
    in_hole_num = 'bx;
    in_hole_suit = 'bx;
    in_pub_num = 'bx;
    in_pub_suit = 'bx;
	
    force clk = 0;
    #CYCLE; rst_n = 0; 
    #CYCLE; rst_n = 1;
    if(out_valid !== 'b0 || out_win_rate !== 'b0) begin //out!==0
        $display("************************************************************");  
        $display("                          FAIL!                              ");    
        $display("*  Output signal should be 0 after initial RESET  at %8t   *",$time);
        $display("************************************************************");
        repeat(2) #CYCLE;
        $finish;
    end
	#CYCLE; release clk;
end endtask


task input_task; begin
	for(j=0; j<9; j=j+1)begin
		$fscanf(file_in, "%d %d %d %d", hcn[j][1], hcs[j][1], hcn[j][0], hcs[j][0]);	
	end	
    $fscanf(file_in, "%d %d %d %d %d %d", pcn[2], pcs[2], pcn[1], pcs[1], pcn[0], pcs[0]);	
    $fscanf(file_in, "%d %d %d %d %d %d %d %d %d", golden_win_rate[0], golden_win_rate[1], golden_win_rate[2], golden_win_rate[3], golden_win_rate[4], golden_win_rate[5], golden_win_rate[6], golden_win_rate[7], golden_win_rate[8]);	
	@(negedge clk);
	in_valid = 'b1;
	in_hole_num  = {hcn[8][1], hcn[8][0], hcn[7][1], hcn[7][0], hcn[6][1], hcn[6][0], hcn[5][1], hcn[5][0], hcn[4][1], hcn[4][0], hcn[3][1], hcn[3][0], hcn[2][1], hcn[2][0], hcn[1][1], hcn[1][0], hcn[0][1], hcn[0][0]};
	in_hole_suit = {hcs[8][1], hcs[8][0], hcs[7][1], hcs[7][0], hcs[6][1], hcs[6][0], hcs[5][1], hcs[5][0], hcs[4][1], hcs[4][0], hcs[3][1], hcs[3][0], hcs[2][1], hcs[2][0], hcs[1][1], hcs[1][0], hcs[0][1], hcs[0][0]};
	in_pub_num = {pcn[2], pcn[1], pcn[0]};
	in_pub_suit = {pcs[2], pcs[1], pcs[0]};
    check_out_valid_task;
	@(negedge clk);

    in_valid = 'b0;
    in_hole_num = 'bx;
    in_hole_suit = 'bx;
    in_pub_num = 'bx;
    in_pub_suit = 'bx;
	@(negedge clk);
end endtask

task wait_out_task; begin
	out_latency = 1;
	while(out_valid !== 1)begin
		if(out_latency === 1001) begin
			$display("********************************************************");     
			$display("*                     FAIL!                            *");
			$display("*  The execution latency are over 1000 cycles          *");//over max
			$display("********************************************************");
			repeat(2) @(negedge clk);
			$finish;
		end
		out_latency = out_latency + 1;
		@(negedge clk);
	end
end endtask

task check_out_valid_task; begin
	if(out_valid !== 0 )begin
		$display("********************************************************");     
		$display("                     FAIL!                              ");
		$display("*  out_valid should not be raised when in_valid is high.  *");
		$display("********************************************************");
		repeat(2) @(negedge clk);
		$finish;
	end
    else if(out_win_rate !== 'b0)begin
		$display("********************************************************");     
		$display("                     FAIL!                              ");
		$display("*  out_win_rate should not be raised when in_valid is high.  *");
		$display("********************************************************");
		repeat(2) @(negedge clk);
		$finish;
	end
end endtask

task check_ans_task; begin
    if(out_win_rate !== golden_out)begin
		$display("[38;2;149;148;154m█[0m[38;2;154;152;158m█[0m[38;2;130;124;130m█[0m[38;2;68;62;64m█[0m[38;2;140;139;142m█[0m[38;2;152;151;156m█[0m[38;2;153;152;157m█[0m[38;2;152;151;156m█[0m[38;2;151;150;155m██[0m[38;2;155;153;158m█[0m[38;2;94;87;89m█[0m[38;2;94;88;92m█[0m[38;2;153;153;158m█[0m[38;2;150;149;154m█[0m[38;2;151;151;156m█[0m[38;2;151;152;156m██[0m[38;2;153;152;158m█[0m[38;2;155;153;158m█[0m[38;2;126;121;125m█[0m[38;2;79;73;76m█[0m[38;2;153;148;155m█[0m[38;2;152;151;157m█[0m[38;2;149;148;154m██[0m[38;2;150;150;155m█[0m[38;2;124;115;120m█[0m[38;2;84;67;69m█[0m[38;2;83;77;78m█[0m[38;2;144;143;147m█[0m[38;2;149;149;155m█[0m[38;2;152;151;157m█[0m[38;2;151;152;156m█[0m[38;2;153;152;158m█[0m[38;2;157;155;161m█[0m[38;2;107;104;105m█[0m[38;2;97;94;96m█[0m[38;2;150;149;154m█[0m[38;2;147;146;152m█[0m[38;2;148;147;153m██[0m[38;2;154;153;159m█[0m[38;2;103;99;104m█[0m[38;2;97;91;96m█[0m[38;2;153;152;157m█[0m[38;2;149;148;154m██[0m[38;2;148;148;153m█[0m[38;2;152;150;157m█[0m[38;2;136;132;136m█[0m[38;2;75;71;69m█[0m[38;2;141;140;143m█[0m[38;2;147;147;152m█[0m[38;2;148;147;153m█[0m[38;2;150;149;155m█[0m[38;2;148;147;151m█[0m[38;2;78;74;75m█[0m[38;2;128;127;130m█[0m[38;2;143;136;139m█[0m[38;2;93;73;72m█[0m[38;2;152;148;150m█[0m[38;2;152;151;156m█[0m[38;2;152;149;154m█[0m[38;2;89;83;85m█[0m[38;2;117;113;116m█[0m[38;2;152;151;155m█[0m[38;2;149;147;152m█[0m[38;2;135;131;137m█[0m[38;2;142;140;145m█[0m[38;2;151;149;156m█[0m[38;2;151;149;155m█[0m[38;2;130;127;130m█[0m[38;2;71;65;68m█[0m[38;2;139;136;141m█[0m[38;2;149;148;153m██[0m[38;2;150;149;155m███[0m[38;2;153;151;157m█[0m[38;2;89;85;88m█[0m[38;2;111;106;110m█[0m[38;2;149;148;154m█[0m[38;2;147;147;153m█[0m[38;2;148;147;153m███[0m[38;2;147;146;152m█[0m[38;2;152;149;155m█[0m[38;2;95;90;95m█[0m[38;2;118;115;119m█[0m[38;2;159;158;163m█[0m[38;2;125;114;117m█[0m[38;2;106;91;95m█[0m[38;2;151;150;154m█[0m[38;2;152;151;157m█[0m[38;2;156;155;160m█[0m[38;2;106;105;105m█[0m[38;2;96;95;96m█[0m");
		$display("[38;2;149;149;155m█[0m[38;2;154;153;159m█[0m[38;2;131;127;131m█[0m[38;2;68;62;63m█[0m[38;2;143;140;145m█[0m[38;2;155;153;159m█[0m[38;2;151;150;155m█[0m[38;2;152;151;156m██[0m[38;2;151;150;156m█[0m[38;2;155;153;157m█[0m[38;2;98;90;96m█[0m[38;2;88;82;86m█[0m[38;2;150;149;154m█[0m[38;2;148;147;153m█[0m[38;2;150;150;156m█[0m[38;2;151;150;156m█[0m[38;2;149;148;154m██[0m[38;2;152;151;157m█[0m[38;2;125;119;123m█[0m[38;2;84;80;80m█[0m[38;2;155;153;159m█[0m[38;2;153;153;159m█[0m[38;2;150;149;155m█[0m[38;2;151;150;156m█[0m[38;2;152;151;157m█[0m[38;2;151;149;154m█[0m[38;2;111;103;105m█[0m[38;2;77;65;68m█[0m[38;2;133;126;129m█[0m[38;2;154;154;158m█[0m[38;2;154;153;159m█[0m[38;2;150;149;155m██[0m[38;2;154;153;158m█[0m[38;2;96;93;95m█[0m[38;2;106;104;105m█[0m[38;2;153;153;158m█[0m[38;2;150;149;155m██[0m[38;2;151;150;155m█[0m[38;2;153;151;156m█[0m[38;2;133;131;136m█[0m[38;2;131;130;135m█[0m[38;2;153;152;157m█[0m[38;2;150;149;155m██[0m[38;2;149;148;154m█[0m[38;2;155;153;159m█[0m[38;2;136;132;136m█[0m[38;2;76;69;72m█[0m[38;2;147;145;149m█[0m[38;2;150;149;155m██[0m[38;2;152;151;157m█[0m[38;2;152;151;156m█[0m[38;2;112;107;111m█[0m[38;2;147;146;150m█[0m[38;2;136;129;132m█[0m[38;2;99;80;80m█[0m[38;2;155;153;157m█[0m[38;2;151;150;156m█[0m[38;2;150;148;153m█[0m[38;2;84;79;80m█[0m[38;2;120;116;119m█[0m[38;2;155;153;159m█[0m[38;2;152;150;155m█[0m[38;2;137;130;137m█[0m[38;2;141;137;143m█[0m[38;2;153;151;158m█[0m[38;2;152;150;156m█[0m[38;2;129;126;130m█[0m[38;2;70;66;68m█[0m[38;2;142;140;144m█[0m[38;2;151;149;155m█[0m[38;2;151;150;156m█[0m[38;2;151;151;156m██[0m[38;2;150;149;154m█[0m[38;2;152;150;155m█[0m[38;2;86;80;84m█[0m[38;2;118;114;117m█[0m[38;2;154;153;159m█[0m[38;2;150;149;155m█[0m[38;2;149;148;154m█[0m[38;2;150;149;155m███[0m[38;2;152;149;156m█[0m[38;2;97;91;96m█[0m[38;2;114;110;114m█[0m[38;2;158;157;162m█[0m[38;2;148;143;145m█[0m[38;2;96;77;80m█[0m[38;2;144;141;146m█[0m[38;2;150;150;156m█[0m[38;2;153;152;158m█[0m[38;2;102;100;101m█[0m[38;2;105;104;105m█[0m");
		$display("[38;2;152;151;157m█[0m[38;2;155;155;161m█[0m[38;2;134;130;134m█[0m[38;2;69;62;64m█[0m[38;2;144;141;146m█[0m[38;2;159;157;164m█[0m[38;2;133;125;132m█[0m[38;2;136;128;133m█[0m[38;2;155;151;156m█[0m[38;2;150;150;155m█[0m[38;2;155;154;158m█[0m[38;2;100;93;98m█[0m[38;2;83;79;82m█[0m[38;2;153;152;157m█[0m[38;2;153;152;158m█[0m[38;2;149;148;154m█[0m[38;2;152;150;156m█[0m[38;2;150;149;155m█[0m[38;2;150;150;156m█[0m[38;2;155;153;159m█[0m[38;2;120;115;118m█[0m[38;2;94;90;91m█[0m[38;2;157;156;162m█[0m[38;2;154;153;159m█[0m[38;2;152;151;157m██[0m[38;2;153;152;158m█[0m[38;2;156;155;161m█[0m[38;2;123;119;122m█[0m[38;2;90;81;80m█[0m[38;2;118;104;104m█[0m[38;2;112;96;98m█[0m[38;2;142;136;139m█[0m[38;2;152;152;156m█[0m[38;2;149;148;155m█[0m[38;2;152;151;156m█[0m[38;2;88;84;87m█[0m[38;2;120;118;119m█[0m[38;2;158;158;162m█[0m[38;2;151;150;155m█[0m[38;2;150;149;153m█[0m[38;2;152;151;155m█[0m[38;2;156;155;160m█[0m[38;2;120;119;123m█[0m[38;2;132;131;136m█[0m[38;2;155;154;160m█[0m[38;2;152;151;156m██[0m[38;2;152;151;157m█[0m[38;2;154;154;159m█[0m[38;2;142;141;144m█[0m[38;2;112;108;112m█[0m[38;2;154;150;157m█[0m[38;2;152;150;156m█[0m[38;2;151;150;156m█[0m[38;2;153;152;157m█[0m[38;2;148;147;153m█[0m[38;2;114;112;118m█[0m[38;2;150;147;154m█[0m[38;2;153;152;156m█[0m[38;2;150;146;150m█[0m[38;2;157;156;161m█[0m[38;2;154;153;158m█[0m[38;2;152;152;157m█[0m[38;2;82;75;77m█[0m[38;2;127;122;126m█[0m[38;2;159;158;164m█[0m[38;2;153;152;159m█[0m[38;2;154;153;159m█[0m[38;2;155;154;160m█[0m[38;2;154;153;159m█[0m[38;2;155;154;159m█[0m[38;2;129;126;130m█[0m[38;2;73;69;70m█[0m[38;2;148;147;152m█[0m[38;2;153;153;158m█[0m[38;2;151;150;155m██[0m[38;2;152;151;157m██[0m[38;2;153;150;156m█[0m[38;2;85;78;82m█[0m[38;2;128;125;129m█[0m[38;2;157;156;162m█[0m[38;2;153;152;158m█[0m[38;2;154;153;159m█[0m[38;2;154;153;158m█[0m[38;2;154;153;159m█[0m[38;2;154;154;160m█[0m[38;2;157;155;160m█[0m[38;2;99;94;97m█[0m[38;2;106;102;104m█[0m[38;2;158;158;162m█[0m[38;2;153;152;153m█[0m[38;2;93;73;71m█[0m[38;2;140;136;140m█[0m[38;2;152;152;158m█[0m[38;2;154;150;156m█[0m[38;2;94;90;92m█[0m[38;2;113;112;112m█[0m");
		$display("[38;2;110;95;97m█[0m[38;2;150;145;149m█[0m[38;2;142;139;142m█[0m[38;2;68;64;64m█[0m[38;2;142;141;146m█[0m[38;2;158;156;162m█[0m[38;2;149;144;150m█[0m[38;2;130;122;127m█[0m[38;2;137;133;137m█[0m[38;2;141;137;143m█[0m[38;2;156;156;158m█[0m[38;2;99;94;98m█[0m[38;2;88;84;88m█[0m[38;2;158;155;161m█[0m[38;2;137;131;139m█[0m[38;2;144;141;148m█[0m[38;2;148;147;153m█[0m[38;2;154;153;159m█[0m[38;2;155;154;160m█[0m[38;2;157;156;162m█[0m[38;2;109;105;109m█[0m[38;2;104;99;101m█[0m[38;2;158;156;162m█[0m[38;2;154;153;160m█[0m[38;2;154;153;159m█[0m[38;2;153;152;158m█[0m[38;2;154;153;159m█[0m[38;2;160;157;164m█[0m[38;2;118;113;116m█[0m[38;2;96;93;91m█[0m[38;2;129;116;115m█[0m[38;2;93;72;69m█[0m[38;2;97;76;73m█[0m[38;2;112;95;98m█[0m[38;2;149;145;149m█[0m[38;2;152;150;153m█[0m[38;2;83;77;78m█[0m[38;2;85;74;74m█[0m[38;2;101;84;84m█[0m[38;2;110;93;93m█[0m[38;2;120;107;106m█[0m[38;2;117;104;104m█[0m[38;2;109;96;96m█[0m[38;2;115;104;106m█[0m[38;2;152;148;152m█[0m[38;2;158;157;163m█[0m[38;2;157;156;162m█[0m[38;2;156;156;162m█[0m[38;2;154;152;158m█[0m[38;2;154;151;157m█[0m[38;2;131;126;130m█[0m[38;2;110;105;109m█[0m[38;2;150;146;152m█[0m[38;2;150;148;153m█[0m[38;2;153;153;159m█[0m[38;2;156;156;162m█[0m[38;2;155;155;160m█[0m[38;2;152;152;157m█[0m[38;2;154;154;158m█[0m[38;2;135;130;133m█[0m[38;2;114;102;103m█[0m[38;2;115;101;102m█[0m[38;2;119;105;107m█[0m[38;2;119;106;109m█[0m[38;2;77;68;69m█[0m[38;2;106;100;102m█[0m[38;2;151;149;153m█[0m[38;2;160;160;165m█[0m[38;2;156;155;161m█[0m[38;2;155;155;161m█[0m[38;2;156;155;161m█[0m[38;2;159;157;163m█[0m[38;2;132;128;132m█[0m[38;2;78;74;75m█[0m[38;2;152;150;155m█[0m[38;2;154;153;159m██[0m[38;2;154;153;158m█[0m[38;2;152;152;157m█[0m[38;2;151;151;157m█[0m[38;2;152;150;153m█[0m[38;2;84;79;81m█[0m[38;2;134;133;136m█[0m[38;2;155;154;160m█[0m[38;2;153;152;158m█[0m[38;2;154;153;159m█[0m[38;2;156;155;161m█[0m[38;2;155;153;159m█[0m[38;2;148;143;149m█[0m[38;2;161;158;163m█[0m[38;2;102;97;100m█[0m[38;2;103;100;103m█[0m[38;2;163;163;166m█[0m[38;2;122;109;112m█[0m[38;2;102;85;87m█[0m[38;2;154;153;157m█[0m[38;2;154;152;159m█[0m[38;2;154;151;154m█[0m[38;2;85;81;82m█[0m[38;2;120;119;120m█[0m");
		$display("[38;2;130;120;122m█[0m[38;2;108;92;93m█[0m[38;2;114;101;101m█[0m[38;2;70;65;65m█[0m[38;2;142;142;147m█[0m[38;2;156;155;161m█[0m[38;2;153;152;158m█[0m[38;2;154;153;159m█[0m[38;2;144;139;146m█[0m[38;2;146;144;150m█[0m[38;2;158;158;161m█[0m[38;2;100;94;98m█[0m[38;2;93;87;92m█[0m[38;2;162;158;164m█[0m[38;2;145;141;148m█[0m[38;2;158;155;162m█[0m[38;2;156;155;161m█[0m[38;2;157;156;161m█[0m[38;2;157;157;163m█[0m[38;2;160;159;165m█[0m[38;2;105;102;107m█[0m[38;2;115;112;115m█[0m[38;2;159;158;163m█[0m[38;2;153;152;158m█[0m[38;2;154;153;159m██[0m[38;2;155;154;160m█[0m[38;2;161;160;167m█[0m[38;2;123;121;123m█[0m[38;2;70;58;58m█[0m[38;2;105;83;83m█[0m[38;2;126;112;110m█[0m[38;2;128;117;119m█[0m[38;2;144;134;136m█[0m[38;2;123;110;111m█[0m[38;2;85;68;68m█[0m[38;2;72;61;60m█[0m[38;2;149;142;139m█[0m[38;2;225;219;216m█[0m[38;2;242;239;237m█[0m[38;2;229;225;224m█[0m[38;2;232;229;226m█[0m[38;2;221;217;214m█[0m[38;2;143;128;126m█[0m[38;2;88;69;67m█[0m[38;2;150;144;147m█[0m[38;2;125;116;118m█[0m[38;2;102;85;86m█[0m[38;2;98;78;76m█[0m[38;2;100;79;76m█[0m[38;2;102;82;80m█[0m[38;2;104;84;82m█[0m[38;2;101;81;79m█[0m[38;2;99;79;77m█[0m[38;2;98;79;78m█[0m[38;2;107;92;92m█[0m[38;2;131;122;126m█[0m[38;2;157;155;159m█[0m[38;2;115;102;105m█[0m[38;2;104;84;85m█[0m[38;2;194;185;182m█[0m[38;2;222;217;213m█[0m[38;2;242;238;235m█[0m[38;2;232;227;225m█[0m[38;2;99;91;91m█[0m[38;2;127;114;115m█[0m[38;2;108;88;90m█[0m[38;2;115;102;105m█[0m[38;2;155;154;159m█[0m[38;2;154;153;159m██[0m[38;2;160;158;163m█[0m[38;2;134;129;133m█[0m[38;2;80;76;77m█[0m[38;2;156;154;158m█[0m[38;2;157;156;161m█[0m[38;2;150;148;154m█[0m[38;2;154;153;159m███[0m[38;2;150;149;152m█[0m[38;2;83;80;83m█[0m[38;2;141;139;142m█[0m[38;2;156;154;160m█[0m[38;2;155;154;160m█[0m[38;2;155;154;159m█[0m[38;2;148;144;149m█[0m[38;2;142;137;142m█[0m[38;2;126;117;122m█[0m[38;2;160;160;164m█[0m[38;2;103;99;99m█[0m[38;2;116;112;115m█[0m[38;2;142;132;135m█[0m[38;2;95;73;74m█[0m[38;2;147;143;145m█[0m[38;2;153;154;159m█[0m[38;2;154;153;158m█[0m[38;2;153;151;155m█[0m[38;2;82;78;78m█[0m[38;2;130;128;132m█[0m");
		$display("[38;2;161;162;166m█[0m[38;2;157;156;160m█[0m[38;2;126;117;120m█[0m[38;2;69;61;60m█[0m[38;2;116;103;107m█[0m[38;2;155;152;157m█[0m[38;2;164;163;169m█[0m[38;2;160;160;166m█[0m[38;2;158;157;163m█[0m[38;2;156;155;161m█[0m[38;2;160;159;163m█[0m[38;2;100;94;97m█[0m[38;2;97;91;95m█[0m[38;2;165;161;167m█[0m[38;2;158;160;164m█[0m[38;2;155;154;160m█[0m[38;2;157;156;161m█[0m[38;2;159;158;163m█[0m[38;2;158;159;163m█[0m[38;2;162;161;167m█[0m[38;2;107;102;108m█[0m[38;2;124;122;124m█[0m[38;2;160;160;165m█[0m[38;2;158;157;163m█[0m[38;2;157;156;162m█[0m[38;2;156;156;162m█[0m[38;2;158;158;164m█[0m[38;2;143;139;142m█[0m[38;2;98;86;87m█[0m[38;2;77;64;64m█[0m[38;2;134;123;123m█[0m[38;2;143;138;140m█[0m[38;2;159;158;163m█[0m[38;2;122;109;113m█[0m[38;2;87;65;66m█[0m[38;2;202;192;190m█[0m[38;2;99;93;90m█[0m[38;2;176;179;181m█[0m[38;2;241;253;255m█[0m[38;2;211;215;218m█[0m[38;2;180;174;172m█[0m[38;2;247;245;244m█[0m[38;2;254;253;254m█[0m[38;2;249;247;246m█[0m[38;2;91;66;63m█[0m[38;2;82;58;57m█[0m[38;2;115;95;93m█[0m[38;2;137;118;116m█[0m[38;2;139;121;117m█[0m[38;2;132;113;111m█[0m[38;2;125;106;104m█[0m[38;2;126;107;104m█[0m[38;2;132;111;110m█[0m[38;2;136;117;115m█[0m[38;2;139;120;117m█[0m[38;2;132;113;110m█[0m[38;2;108;87;84m█[0m[38;2;93;72;72m█[0m[38;2;70;44;44m█[0m[38;2;207;198;194m█[0m[38;2;255;255;255m█[0m[38;2;181;174;174m█[0m[38;2;216;213;212m█[0m[38;2;240;244;244m█[0m[38;2;89;86;85m█[0m[38;2;205;202;201m█[0m[38;2;241;237;236m█[0m[38;2;126;109;109m█[0m[38;2;97;83;84m█[0m[38;2;158;156;161m█[0m[38;2;156;155;161m█[0m[38;2;157;156;161m█[0m[38;2;135;132;135m█[0m[38;2;90;86;87m█[0m[38;2;150;147;149m█[0m[38;2;148;145;148m█[0m[38;2;135;131;136m█[0m[38;2;152;151;156m█[0m[38;2;158;157;162m██[0m[38;2;148;147;150m█[0m[38;2;82;80;82m█[0m[38;2;149;147;150m█[0m[38;2;157;156;162m█[0m[38;2;156;155;161m█[0m[38;2;156;155;159m█[0m[38;2;129;122;125m█[0m[38;2;139;135;137m█[0m[38;2;151;150;153m█[0m[38;2;163;162;167m█[0m[38;2;107;103;105m█[0m[38;2;97;88;88m█[0m[38;2;102;80;83m█[0m[38;2;143;134;137m█[0m[38;2;158;159;162m█[0m[38;2;156;155;160m█[0m[38;2;157;156;161m█[0m[38;2;154;151;155m█[0m[38;2;81;77;78m█[0m[38;2;135;133;137m█[0m");
		$display("[38;2;159;159;164m██[0m[38;2;148;145;151m█[0m[38;2;76;68;70m█[0m[38;2;116;103;102m█[0m[38;2;107;88;87m█[0m[38;2;129;115;117m█[0m[38;2;156;153;157m█[0m[38;2;160;160;164m█[0m[38;2;157;157;163m█[0m[38;2;162;160;165m█[0m[38;2;100;94;97m█[0m[38;2;100;95;99m█[0m[38;2;166;163;169m█[0m[38;2;160;160;166m█[0m[38;2;161;160;166m███[0m[38;2;160;160;165m█[0m[38;2;165;164;169m█[0m[38;2;108;105;109m█[0m[38;2;128;127;129m█[0m[38;2;167;167;172m█[0m[38;2;164;164;170m█[0m[38;2;163;162;168m█[0m[38;2;153;147;153m█[0m[38;2;127;115;118m█[0m[38;2;122;109;110m█[0m[38;2;114;104;106m█[0m[38;2;84;79;82m█[0m[38;2;163;160;165m█[0m[38;2;164;163;169m█[0m[38;2;154;150;155m█[0m[38;2;76;55;53m█[0m[38;2;209;200;199m█[0m[38;2;253;255;255m█[0m[38;2;100;96;97m█[0m[38;2;146;162;169m█[0m[38;2;205;236;248m█[0m[38;2;145;147;154m█[0m[38;2;236;232;231m█[0m[38;2;251;250;250m█[0m[38;2;252;251;252m█[0m[38;2;226;221;221m█[0m[38;2;73;46;46m█[0m[38;2;82;57;55m█[0m[38;2;103;82;79m█[0m[38;2;110;88;86m█[0m[38;2;125;105;103m█[0m[38;2;140;121;120m█[0m[38;2;150;132;132m█[0m[38;2;150;132;131m█[0m[38;2;146;125;126m█[0m[38;2;134;114;115m█[0m[38;2;118;97;97m█[0m[38;2;103;80;80m█[0m[38;2;96;72;72m█[0m[38;2;68;38;40m█[0m[38;2;61;32;34m█[0m[38;2;206;198;195m█[0m[38;2;255;255;255m█[0m[38;2;218;210;210m█[0m[38;2;127;125;128m█[0m[38;2;203;230;240m█[0m[38;2;81;82;81m█[0m[38;2;176;190;196m█[0m[38;2;245;252;255m█[0m[38;2;248;244;243m█[0m[38;2;92;71;70m█[0m[38;2;130;121;125m█[0m[38;2;161;161;167m█[0m[38;2;161;159;165m█[0m[38;2;139;135;140m█[0m[38;2;101;96;99m█[0m[38;2;149;145;149m█[0m[38;2;144;141;146m█[0m[38;2;161;161;166m█[0m[38;2;159;158;164m██[0m[38;2;162;161;167m█[0m[38;2;148;147;150m█[0m[38;2;83;80;82m█[0m[38;2;156;154;158m█[0m[38;2;158;157;162m█[0m[38;2;158;157;163m█[0m[38;2;161;160;166m█[0m[38;2;160;160;165m█[0m[38;2;160;160;164m█[0m[38;2;161;160;166m█[0m[38;2;167;167;172m█[0m[38;2;110;104;106m█[0m[38;2;83;69;71m█[0m[38;2;148;138;142m█[0m[38;2;161;159;165m█[0m[38;2;157;157;162m█[0m[38;2;159;158;163m██[0m[38;2;156;154;158m█[0m[38;2;82;78;78m█[0m[38;2;140;138;142m█[0m");
		$display("[38;2;162;161;167m█[0m[38;2;160;160;166m█[0m[38;2;149;146;150m█[0m[38;2;80;73;76m█[0m[38;2;154;155;157m█[0m[38;2;158;155;157m█[0m[38;2;124;111;112m█[0m[38;2;104;87;86m█[0m[38;2;124;112;112m█[0m[38;2;152;148;151m█[0m[38;2;167;164;169m█[0m[38;2;99;94;98m█[0m[38;2;101;98;102m█[0m[38;2;169;168;173m█[0m[38;2;164;165;171m█[0m[38;2;165;165;171m█[0m[38;2;165;164;170m█[0m[38;2;162;161;166m█[0m[38;2;158;156;162m█[0m[38;2;158;154;159m█[0m[38;2;108;103;103m█[0m[38;2;108;101;101m█[0m[38;2;141;132;134m█[0m[38;2;133;120;122m█[0m[38;2;130;119;121m█[0m[38;2;134;123;126m█[0m[38;2;146;139;143m█[0m[38;2;166;165;169m█[0m[38;2;120;117;120m█[0m[38;2;89;85;89m█[0m[38;2;166;165;170m█[0m[38;2;164;163;169m█[0m[38;2;151;144;150m█[0m[38;2;84;64;63m█[0m[38;2;242;238;236m█[0m[38;2;232;246;249m█[0m[38;2;107;111;114m█[0m[38;2;128;135;136m█[0m[38;2;161;173;180m█[0m[38;2;114;105;109m█[0m[38;2;229;223;221m█[0m[38;2;252;250;251m█[0m[38;2;255;255;255m█[0m[38;2;168;155;154m█[0m[38;2;55;27;26m█[0m[38;2;151;133;131m█[0m[38;2;172;159;156m█[0m[38;2;157;142;139m█[0m[38;2;140;121;118m█[0m[38;2;124;105;102m█[0m[38;2;117;98;96m█[0m[38;2;118;99;96m█[0m[38;2;126;105;103m█[0m[38;2;135;114;113m█[0m[38;2;146;129;127m█[0m[38;2;160;146;142m█[0m[38;2;167;155;152m█[0m[38;2;115;94;92m█[0m[38;2;66;37;38m█[0m[38;2;222;217;214m█[0m[38;2;255;255;255m█[0m[38;2;185;175;174m█[0m[38;2;99;91;93m█[0m[38;2;162;177;182m█[0m[38;2;80;79;78m█[0m[38;2;173;193;204m█[0m[38;2;220;240;245m█[0m[38;2;255;255;254m█[0m[38;2;111;91;87m█[0m[38;2;118;107;109m█[0m[38;2;164;164;170m█[0m[38;2;162;161;167m█[0m[38;2;134;132;136m█[0m[38;2;104;101;104m█[0m[38;2;167;165;172m█[0m[38;2;164;162;168m█[0m[38;2;162;161;167m█[0m[38;2;160;159;165m█[0m[38;2;159;158;164m█[0m[38;2;162;161;167m█[0m[38;2;146;144;146m█[0m[38;2;82;79;79m█[0m[38;2;157;154;159m█[0m[38;2;160;159;165m█[0m[38;2;160;159;166m█[0m[38;2;161;160;166m█[0m[38;2;162;161;167m█[0m[38;2;163;163;169m█[0m[38;2;165;165;171m█[0m[38;2;136;125;129m█[0m[38;2;82;68;72m█[0m[38;2;123;120;123m█[0m[38;2;166;165;171m█[0m[38;2;161;160;166m█[0m[38;2;162;161;167m██[0m[38;2;163;162;167m█[0m[38;2;157;155;159m█[0m[38;2;80;76;77m█[0m[38;2;142;139;144m█[0m");
		$display("[38;2;162;161;167m█[0m[38;2;164;163;169m█[0m[38;2;154;152;155m█[0m[38;2;83;77;77m█[0m[38;2;154;154;157m█[0m[38;2;165;166;171m█[0m[38;2;165;165;169m█[0m[38;2;156;153;155m█[0m[38;2;130;117;119m█[0m[38;2;111;95;96m█[0m[38;2;120;105;107m█[0m[38;2;89;79;81m█[0m[38;2;94;85;87m█[0m[38;2;136;126;128m█[0m[38;2;132;119;122m█[0m[38;2;127;114;115m█[0m[38;2;122;108;110m█[0m[38;2;120;105;107m██[0m[38;2;125;109;112m█[0m[38;2;102;91;94m█[0m[38;2;86;77;77m█[0m[38;2;140;130;132m█[0m[38;2;146;140;143m█[0m[38;2;157;154;158m█[0m[38;2;165;162;169m█[0m[38;2;165;163;170m█[0m[38;2;168;168;173m█[0m[38;2;115;113;117m█[0m[38;2;103;100;104m█[0m[38;2;169;169;173m█[0m[38;2;165;165;170m█[0m[38;2;167;165;170m█[0m[38;2;101;86;85m█[0m[38;2;166;153;150m█[0m[38;2;253;255;255m█[0m[38;2;136;140;141m█[0m[38;2;140;154;161m█[0m[38;2;181;200;206m█[0m[38;2;136;133;136m█[0m[38;2;196;186;186m█[0m[38;2;254;253;253m██[0m[38;2;187;178;179m█[0m[38;2;78;54;52m█[0m[38;2;109;87;84m█[0m[38;2;120;102;98m█[0m[38;2;136;119;117m█[0m[38;2;153;136;135m█[0m[38;2;165;151;149m█[0m[38;2;171;157;158m██[0m[38;2;166;151;151m█[0m[38;2;154;140;138m█[0m[38;2;141;123;122m█[0m[38;2;124;104;102m█[0m[38;2;114;94;92m█[0m[38;2;111;92;90m█[0m[38;2;174;163;162m█[0m[38;2;252;252;251m█[0m[38;2;239;236;235m█[0m[38;2;121;106;106m█[0m[38;2;140;142;143m█[0m[38;2;175;192;196m█[0m[38;2;90;89;92m█[0m[38;2;180;200;208m█[0m[38;2;240;254;255m█[0m[38;2;220;215;213m█[0m[38;2;77;49;47m█[0m[38;2;106;89;90m█[0m[38;2;159;157;161m█[0m[38;2;163;160;164m█[0m[38;2;129;124;127m█[0m[38;2;109;104;107m█[0m[38;2;169;168;173m█[0m[38;2;165;164;170m█[0m[38;2;164;164;170m█[0m[38;2;163;162;168m█[0m[38;2;159;158;164m█[0m[38;2;162;161;167m█[0m[38;2;144;143;145m█[0m[38;2;82;77;77m█[0m[38;2;158;157;162m█[0m[38;2;162;163;169m█[0m[38;2;163;161;168m█[0m[38;2;163;161;167m█[0m[38;2;160;159;163m█[0m[38;2;152;148;151m█[0m[38;2;122;105;106m█[0m[38;2;116;98;100m█[0m[38;2;104;98;99m█[0m[38;2;124;121;123m█[0m[38;2;166;165;170m█[0m[38;2;162;161;167m██[0m[38;2;163;162;168m█[0m[38;2;165;164;170m█[0m[38;2;160;158;161m█[0m[38;2;81;77;78m█[0m[38;2;142;139;143m█[0m");
		$display("[38;2;161;160;166m█[0m[38;2;163;162;167m█[0m[38;2;152;149;153m█[0m[38;2;76;70;72m█[0m[38;2;150;150;154m█[0m[38;2;167;167;172m█[0m[38;2;165;164;170m█[0m[38;2;165;165;171m█[0m[38;2;168;167;173m█[0m[38;2;164;162;167m█[0m[38;2;156;151;155m█[0m[38;2;100;92;94m█[0m[38;2;83;67;66m█[0m[38;2;111;92;92m█[0m[38;2;148;142;142m█[0m[38;2;150;145;148m█[0m[38;2;155;149;154m█[0m[38;2;157;155;160m█[0m[38;2;161;160;166m█[0m[38;2;167;167;172m█[0m[38;2;129;125;128m█[0m[38;2;91;86;87m█[0m[38;2;169;168;174m█[0m[38;2;163;163;169m█[0m[38;2;162;161;167m██[0m[38;2;164;163;169m█[0m[38;2;169;168;173m█[0m[38;2;101;100;102m█[0m[38;2;109;108;109m█[0m[38;2;170;169;174m█[0m[38;2;167;166;171m██[0m[38;2;161;159;163m█[0m[38;2;108;93;95m█[0m[38;2;150;138;136m█[0m[38;2;149;141;142m█[0m[38;2;147;146;149m█[0m[38;2;226;222;222m█[0m[38;2;245;243;242m█[0m[38;2;250;249;249m█[0m[38;2;250;247;248m█[0m[38;2;249;247;248m█[0m[38;2;252;249;250m█[0m[38;2;236;233;232m█[0m[38;2;244;241;240m█[0m[38;2;253;252;251m█[0m[38;2;255;255;255m████████[0m[38;2;255;254;254m█[0m[38;2;249;248;248m█[0m[38;2;245;243;245m█[0m[38;2;254;253;254m█[0m[38;2;249;247;248m█[0m[38;2;249;246;247m█[0m[38;2;246;243;244m█[0m[38;2;230;226;226m█[0m[38;2;199;196;195m█[0m[38;2;98;95;95m█[0m[38;2;212;213;213m█[0m[38;2;203;194;193m█[0m[38;2;104;89;88m█[0m[38;2;141;151;162m█[0m[38;2;119;122;129m█[0m[38;2;116;112;114m█[0m[38;2;181;206;218m█[0m[38;2;121;127;131m█[0m[38;2;116;114;118m█[0m[38;2;170;172;179m█[0m[38;2;168;167;172m█[0m[38;2;162;159;163m█[0m[38;2;156;151;156m█[0m[38;2;161;159;164m█[0m[38;2;169;168;174m█[0m[38;2;144;141;143m█[0m[38;2;77;71;72m█[0m[38;2;131;119;121m█[0m[38;2;127;113;115m█[0m[38;2;123;109;110m█[0m[38;2;118;101;100m█[0m[38;2;117;97;96m█[0m[38;2;97;72;70m█[0m[38;2;114;92;92m█[0m[38;2;156;146;149m█[0m[38;2;116;112;116m█[0m[38;2;125;120;124m█[0m[38;2;168;167;173m█[0m[38;2;162;161;167m█[0m[38;2;161;160;166m█[0m[38;2;162;161;167m█[0m[38;2;164;163;169m█[0m[38;2;161;160;162m█[0m[38;2;81;78;79m█[0m[38;2;140;139;142m█[0m");
		$display("[38;2;161;160;166m█[0m[38;2;163;162;168m█[0m[38;2;156;154;159m█[0m[38;2;77;70;74m█[0m[38;2;143;141;146m█[0m[38;2;168;167;173m█[0m[38;2;167;166;172m████[0m[38;2;172;171;175m█[0m[38;2;106;101;104m█[0m[38;2;73;57;57m█[0m[38;2;154;145;149m█[0m[38;2;171;171;175m█[0m[38;2;168;168;174m█[0m[38;2;167;167;173m█[0m[38;2;166;165;172m█[0m[38;2;166;165;171m█[0m[38;2;170;169;175m█[0m[38;2;118;113;116m█[0m[38;2;95;90;93m█[0m[38;2;171;167;174m█[0m[38;2;166;164;170m█[0m[38;2;165;164;170m█[0m[38;2;164;163;169m█[0m[38;2;165;164;170m█[0m[38;2;167;166;171m█[0m[38;2;93;90;91m█[0m[38;2;113;108;111m█[0m[38;2;169;166;171m█[0m[38;2;167;166;172m█[0m[38;2;166;165;171m█[0m[38;2;171;171;176m█[0m[38;2;167;165;170m█[0m[38;2;113;98;101m█[0m[38;2;82;65;67m█[0m[38;2;155;149;150m█[0m[38;2;255;255;255m█[0m[38;2;250;248;249m█[0m[38;2;249;247;248m████[0m[38;2;251;250;251m█[0m[38;2;250;248;250m█[0m[38;2;249;247;248m██████████[0m[38;2;250;248;249m██[0m[38;2;249;247;248m███[0m[38;2;250;248;249m█[0m[38;2;253;251;252m█[0m[38;2;247;245;245m█[0m[38;2;106;100;99m█[0m[38;2;159;152;151m█[0m[38;2;138;148;154m█[0m[38;2;164;201;216m█[0m[38;2;189;239;255m█[0m[38;2;164;197;212m█[0m[38;2;107;112;119m█[0m[38;2;187;233;251m█[0m[38;2;110;122;130m█[0m[38;2;137;160;170m█[0m[38;2;159;185;194m█[0m[38;2;112;104;108m█[0m[38;2;114;107;108m█[0m[38;2;128;118;121m█[0m[38;2;154;149;152m█[0m[38;2;129;114;115m█[0m[38;2;106;91;90m█[0m[38;2;74;67;65m█[0m[38;2;134;123;126m█[0m[38;2;154;146;150m█[0m[38;2;155;150;151m█[0m[38;2;138;127;128m█[0m[38;2;137;124;125m█[0m[38;2;128;111;111m█[0m[38;2;111;87;88m█[0m[38;2;132;117;120m█[0m[38;2;114;111;115m█[0m[38;2;128;124;127m█[0m[38;2;171;170;175m█[0m[38;2;163;162;168m█[0m[38;2;162;161;167m█[0m[38;2;163;162;168m█[0m[38;2;164;163;169m█[0m[38;2;162;158;162m█[0m[38;2;81;77;79m█[0m[38;2;138;136;141m█[0m");
		$display("[38;2;164;163;169m█[0m[38;2;168;167;173m█[0m[38;2;162;159;165m█[0m[38;2;74;68;73m█[0m[38;2;140;140;143m█[0m[38;2;171;170;175m█[0m[38;2;166;165;170m█[0m[38;2;165;164;170m██[0m[38;2;167;166;172m█[0m[38;2;173;170;174m█[0m[38;2;104;98;101m█[0m[38;2;89;77;79m█[0m[38;2;171;168;173m█[0m[38;2;169;169;174m█[0m[38;2;169;168;174m█[0m[38;2;167;166;172m███[0m[38;2;171;170;174m█[0m[38;2;102;98;99m█[0m[38;2;110;104;107m█[0m[38;2;172;168;174m█[0m[38;2;168;166;171m█[0m[38;2;168;167;173m█[0m[38;2;167;166;172m██[0m[38;2;171;169;174m█[0m[38;2;96;92;95m█[0m[38;2;119;114;119m█[0m[38;2;173;170;177m█[0m[38;2;168;167;173m█[0m[38;2;172;172;176m█[0m[38;2;137;128;130m█[0m[38;2;83;62;64m█[0m[38;2;144;131;130m█[0m[38;2;183;176;174m█[0m[38;2;138;133;133m█[0m[38;2;255;254;254m█[0m[38;2;249;247;248m███████████████████████[0m[38;2;251;249;250m█[0m[38;2;239;237;237m█[0m[38;2;101;99;97m█[0m[38;2;230;229;228m█[0m[38;2;231;235;239m█[0m[38;2;122;121;128m█[0m[38;2;146;173;185m█[0m[38;2;181;228;246m█[0m[38;2;174;216;233m█[0m[38;2;183;226;245m█[0m[38;2;100;110;115m█[0m[38;2;144;166;181m█[0m[38;2;123;135;145m█[0m[38;2;160;193;206m█[0m[38;2;179;221;240m█[0m[38;2;176;201;212m█[0m[38;2;163;166;171m█[0m[38;2;153;148;152m█[0m[38;2;151;144;147m█[0m[38;2;79;75;75m█[0m[38;2;163;162;166m█[0m[38;2;170;170;175m█[0m[38;2;170;169;174m█[0m[38;2;168;166;172m█[0m[38;2;152;143;148m█[0m[38;2;143;133;135m█[0m[38;2;144;132;132m█[0m[38;2;110;87;89m█[0m[38;2;91;81;81m█[0m[38;2;130;129;131m█[0m[38;2;169;168;173m█[0m[38;2;164;164;169m█[0m[38;2;166;165;171m███[0m[38;2;162;159;165m█[0m[38;2;82;77;81m█[0m[38;2;139;137;143m█[0m");
		$display("[38;2;164;163;169m█[0m[38;2;170;168;175m█[0m[38;2;150;149;152m█[0m[38;2;66;65;65m█[0m[38;2;150;149;153m█[0m[38;2;170;169;175m█[0m[38;2;166;165;170m█[0m[38;2;164;163;169m█[0m[38;2;165;164;170m█[0m[38;2;168;167;173m█[0m[38;2;174;172;177m█[0m[38;2;100;92;95m█[0m[38;2;114;108;111m█[0m[38;2;173;172;177m█[0m[38;2;168;167;173m█[0m[38;2;167;166;172m█[0m[38;2;166;165;171m█[0m[38;2;167;166;171m█[0m[38;2;167;166;172m█[0m[38;2;169;168;172m█[0m[38;2;91;87;87m█[0m[38;2;123;118;121m█[0m[38;2;170;167;172m█[0m[38;2;156;153;158m█[0m[38;2;162;159;164m█[0m[38;2;167;166;172m█[0m[38;2;169;168;174m█[0m[38;2;173;171;177m█[0m[38;2;104;99;104m█[0m[38;2;123;119;124m█[0m[38;2;175;173;180m█[0m[38;2;173;172;176m█[0m[38;2;115;101;101m█[0m[38;2;71;45;44m█[0m[38;2;183;172;169m█[0m[38;2;255;255;255m█[0m[38;2;208;205;203m█[0m[38;2;124;122;122m█[0m[38;2;254;252;253m█[0m[38;2;249;247;248m███████████████████████[0m[38;2;252;250;251m█[0m[38;2;230;228;228m█[0m[38;2;95;92;90m█[0m[38;2;232;230;230m█[0m[38;2;255;253;253m█[0m[38;2;216;208;206m█[0m[38;2;86;67;65m█[0m[38;2;129;144;153m█[0m[38;2;186;231;252m█[0m[38;2;179;224;242m█[0m[38;2;96;105;111m█[0m[38;2;159;190;205m█[0m[38;2;183;229;247m█[0m[38;2;181;228;246m█[0m[38;2;176;220;238m█[0m[38;2;160;194;209m█[0m[38;2;146;157;166m█[0m[38;2;140;134;136m█[0m[38;2;140;134;137m█[0m[38;2;79;75;77m█[0m[38;2;161;160;164m█[0m[38;2;171;171;175m█[0m[38;2;169;168;174m██[0m[38;2;170;169;174m█[0m[38;2;164;161;166m█[0m[38;2;165;161;166m█[0m[38;2;150;142;143m█[0m[38;2;84;72;73m█[0m[38;2;133;131;134m█[0m[38;2;172;171;176m█[0m[38;2;165;164;169m█[0m[38;2;165;164;170m█[0m[38;2;166;165;171m█[0m[38;2;168;167;173m█[0m[38;2;167;164;170m█[0m[38;2;83;78;82m█[0m[38;2;138;136;141m█[0m");
		$display("[38;2;166;165;171m█[0m[38;2;171;170;176m█[0m[38;2;139;136;139m█[0m[38;2;69;66;65m█[0m[38;2;158;156;161m█[0m[38;2;168;167;174m█[0m[38;2;167;166;172m██[0m[38;2;169;168;174m█[0m[38;2;172;171;176m█[0m[38;2;173;170;175m█[0m[38;2;93;86;88m█[0m[38;2;120;116;120m█[0m[38;2;172;171;176m█[0m[38;2;167;166;173m█[0m[38;2;167;166;172m███[0m[38;2;168;167;173m█[0m[38;2;170;167;172m█[0m[38;2;86;81;82m█[0m[38;2;130;127;129m█[0m[38;2;165;160;165m█[0m[38;2;143;132;137m█[0m[38;2;148;140;144m█[0m[38;2;168;166;171m█[0m[38;2;172;171;176m█[0m[38;2;176;175;180m█[0m[38;2;112;109;112m█[0m[38;2;121;119;122m█[0m[38;2;177;177;182m█[0m[38;2;128;117;118m█[0m[38;2;66;37;36m█[0m[38;2;198;188;187m█[0m[38;2;255;255;255m█[0m[38;2;255;253;253m█[0m[38;2;211;208;206m█[0m[38;2;118;114;115m█[0m[38;2;253;250;251m█[0m[38;2;249;247;248m███████████████████████[0m[38;2;253;251;252m█[0m[38;2;221;218;218m█[0m[38;2;92;88;87m█[0m[38;2;237;235;235m█[0m[38;2;251;249;250m█[0m[38;2;255;255;255m█[0m[38;2;208;201;199m█[0m[38;2;69;47;47m█[0m[38;2;157;182;196m█[0m[38;2;182;225;243m█[0m[38;2;92;99;104m█[0m[38;2;162;193;208m█[0m[38;2;181;227;246m█[0m[38;2;177;222;240m█[0m[38;2;137;159;173m█[0m[38;2;132;145;157m█[0m[38;2;144;166;180m█[0m[38;2;149;164;172m█[0m[38;2;137;136;138m█[0m[38;2;78;73;75m█[0m[38;2;163;158;162m█[0m[38;2;173;171;176m█[0m[38;2;171;170;176m███[0m[38;2;166;165;171m█[0m[38;2;166;164;170m█[0m[38;2;171;168;174m█[0m[38;2;102;99;100m█[0m[38;2;93;81;83m█[0m[38;2;166;163;166m█[0m[38;2;169;169;174m█[0m[38;2;167;167;172m█[0m[38;2;168;167;173m█[0m[38;2;169;168;174m█[0m[38;2;169;167;171m█[0m[38;2;84;80;81m█[0m[38;2;132;131;135m█[0m");
		$display("[38;2;171;170;176m█[0m[38;2;175;174;179m█[0m[38;2;132;129;131m█[0m[38;2;69;67;66m█[0m[38;2;162;161;165m█[0m[38;2;169;169;173m█[0m[38;2;169;168;174m█[0m[38;2;170;169;175m█[0m[38;2;172;171;177m█[0m[38;2;173;173;178m█[0m[38;2;170;169;173m█[0m[38;2;81;77;76m█[0m[38;2;117;115;118m█[0m[38;2;172;171;177m█[0m[38;2;169;168;174m█[0m[38;2;172;171;177m█[0m[38;2;171;170;176m█[0m[38;2;169;168;174m██[0m[38;2;169;167;172m█[0m[38;2;87;82;84m█[0m[38;2;127;124;125m█[0m[38;2;174;173;178m█[0m[38;2;171;169;174m█[0m[38;2;172;171;176m█[0m[38;2;171;170;176m█[0m[38;2;171;169;175m█[0m[38;2;172;171;177m█[0m[38;2;116;113;116m█[0m[38;2;119;116;119m█[0m[38;2;168;164;168m█[0m[38;2;69;47;46m█[0m[38;2;164;149;146m█[0m[38;2;255;255;255m█[0m[38;2;249;247;248m█[0m[38;2;253;252;252m█[0m[38;2;211;210;208m█[0m[38;2;117;113;113m█[0m[38;2;252;249;250m█[0m[38;2;253;252;253m█[0m[38;2;255;254;254m█[0m[38;2;251;249;250m█[0m[38;2;248;246;246m█[0m[38;2;250;247;248m█[0m[38;2;255;254;254m█[0m[38;2;255;253;254m█[0m[38;2;251;249;250m██[0m[38;2;249;247;248m█[0m[38;2;250;247;248m█[0m[38;2;250;248;249m██[0m[38;2;249;247;248m█[0m[38;2;252;250;251m█[0m[38;2;251;249;250m█[0m[38;2;254;252;254m█[0m[38;2;255;254;255m█[0m[38;2;253;251;252m█[0m[38;2;253;250;251m█[0m[38;2;254;252;253m█[0m[38;2;255;255;255m█[0m[38;2;254;252;253m██[0m[38;2;209;206;207m█[0m[38;2;94;90;89m█[0m[38;2;243;240;241m█[0m[38;2;250;248;249m█[0m[38;2;249;247;248m█[0m[38;2;255;255;255m█[0m[38;2;134;116;115m█[0m[38;2;98;100;108m█[0m[38;2;180;221;239m█[0m[38;2;85;92;93m█[0m[38;2;163;198;213m█[0m[38;2;180;227;245m█[0m[38;2;178;223;243m██[0m[38;2;182;230;246m█[0m[38;2;177;221;239m█[0m[38;2;177;218;236m█[0m[38;2;156;170;177m█[0m[38;2;76;69;72m█[0m[38;2;163;159;163m█[0m[38;2;174;173;178m█[0m[38;2;172;171;176m█[0m[38;2;171;170;176m█[0m[38;2;169;168;174m█[0m[38;2;168;167;173m██[0m[38;2;174;171;176m█[0m[38;2;99;94;96m█[0m[38;2;104;92;92m█[0m[38;2;119;102;102m█[0m[38;2;147;137;138m█[0m[38;2;162;158;162m█[0m[38;2;168;166;171m█[0m[38;2;169;168;173m█[0m[38;2;169;167;171m█[0m[38;2;82;77;78m█[0m[38;2;133;131;134m█[0m");
		$display("[38;2;173;173;178m█[0m[38;2;178;178;182m█[0m[38;2;126;123;125m█[0m[38;2;72;67;68m█[0m[38;2;169;168;173m█[0m[38;2;175;174;179m█[0m[38;2;172;172;177m█[0m[38;2;173;172;178m█[0m[38;2;174;173;179m█[0m[38;2;173;173;179m█[0m[38;2;165;164;168m█[0m[38;2;73;67;67m█[0m[38;2;115;112;115m█[0m[38;2;174;173;179m█[0m[38;2;170;169;175m█[0m[38;2;173;172;178m█[0m[38;2;171;170;176m█[0m[38;2;169;168;174m█[0m[38;2;170;169;175m█[0m[38;2;174;173;177m█[0m[38;2;94;89;91m█[0m[38;2;118;115;117m█[0m[38;2;175;175;180m█[0m[38;2;171;170;176m██[0m[38;2;170;169;175m█[0m[38;2;169;168;174m█[0m[38;2;176;176;182m█[0m[38;2;124;122;123m█[0m[38;2;117;114;116m█[0m[38;2;180;174;177m█[0m[38;2;93;74;71m█[0m[38;2;240;235;234m█[0m[38;2;251;249;249m█[0m[38;2;249;247;248m█[0m[38;2;254;252;252m█[0m[38;2;209;206;205m█[0m[38;2;120;115;114m█[0m[38;2;254;252;252m█[0m[38;2;216;211;210m█[0m[38;2;172;163;163m█[0m[38;2;164;153;153m█[0m[38;2;166;157;156m█[0m[38;2;157;146;145m█[0m[38;2;157;142;142m█[0m[38;2;202;194;194m█[0m[38;2;208;202;203m█[0m[38;2;223;217;219m█[0m[38;2;253;251;252m█[0m[38;2;244;245;246m█[0m[38;2;238;242;243m█[0m[38;2;239;242;243m█[0m[38;2;251;251;252m█[0m[38;2;208;204;204m█[0m[38;2;206;202;202m█[0m[38;2;210;203;203m█[0m[38;2;164;153;153m█[0m[38;2;156;143;142m█[0m[38;2;155;142;138m█[0m[38;2;150;136;134m█[0m[38;2;164;150;150m█[0m[38;2;210;204;204m█[0m[38;2;254;252;253m█[0m[38;2;198;195;196m█[0m[38;2;93;88;87m█[0m[38;2;246;242;243m█[0m[38;2;251;248;249m█[0m[38;2;249;247;248m█[0m[38;2;253;252;252m█[0m[38;2;215;210;210m█[0m[38;2;146;142;147m█[0m[38;2;184;207;215m█[0m[38;2;80;84;85m█[0m[38;2;158;195;211m█[0m[38;2;179;225;244m█[0m[38;2;178;223;242m█[0m[38;2;179;225;243m█[0m[38;2;143;170;182m█[0m[38;2;119;130;138m█[0m[38;2;120;129;139m█[0m[38;2;113;115;120m█[0m[38;2;74;65;68m█[0m[38;2;156;152;156m█[0m[38;2;174;174;178m█[0m[38;2;171;171;176m█[0m[38;2;169;168;174m██[0m[38;2;172;171;177m█[0m[38;2;174;173;179m█[0m[38;2;176;174;179m█[0m[38;2;93;87;89m█[0m[38;2;141;139;141m█[0m[38;2;167;163;168m█[0m[38;2;141;127;131m█[0m[38;2;131;115;117m█[0m[38;2;129;113;114m█[0m[38;2;128;112;112m█[0m[38;2;129;113;114m█[0m[38;2;77;69;68m█[0m[38;2;113;104;104m█[0m");
		$display("[38;2;173;174;179m█[0m[38;2;179;179;183m█[0m[38;2;116;113;116m█[0m[38;2;75;67;70m█[0m[38;2;172;170;174m█[0m[38;2;176;176;181m█[0m[38;2;174;173;179m█[0m[38;2;175;174;180m█[0m[38;2;176;175;181m█[0m[38;2;180;180;185m█[0m[38;2;153;147;152m█[0m[38;2;66;56;59m█[0m[38;2;117;115;118m█[0m[38;2;178;177;182m█[0m[38;2;173;172;178m█[0m[38;2;176;175;181m█[0m[38;2;175;174;180m█[0m[38;2;172;171;177m█[0m[38;2;171;170;176m█[0m[38;2;174;173;177m█[0m[38;2;98;94;96m█[0m[38;2;107;104;107m█[0m[38;2;175;174;180m█[0m[38;2;172;171;177m█[0m[38;2;172;173;178m█[0m[38;2;175;175;180m█[0m[38;2;169;166;171m█[0m[38;2;155;147;149m█[0m[38;2;118;109;109m█[0m[38;2;105;95;95m█[0m[38;2;193;187;187m█[0m[38;2;213;209;208m█[0m[38;2;251;249;249m█[0m[38;2;249;247;248m██[0m[38;2;255;255;254m█[0m[38;2;202;199;198m█[0m[38;2;128;123;123m█[0m[38;2;186;179;177m█[0m[38;2;72;51;51m█[0m[38;2;179;171;169m█[0m[38;2;217;217;216m█[0m[38;2;222;222;220m█[0m[38;2;219;216;214m█[0m[38;2;176;166;164m█[0m[38;2;63;39;37m█[0m[38;2;165;154;152m█[0m[38;2;247;246;246m█[0m[38;2;229;237;240m█[0m[38;2;191;215;219m█[0m[38;2;171;191;198m█[0m[38;2;173;192;200m█[0m[38;2;212;231;237m█[0m[38;2;239;238;238m█[0m[38;2;156;143;140m█[0m[38;2;66;41;39m█[0m[38;2;179;168;166m█[0m[38;2;222;218;218m█[0m[38;2;225;223;220m█[0m[38;2;210;207;203m█[0m[38;2;147;134;132m█[0m[38;2;54;32;31m█[0m[38;2;183;174;172m█[0m[38;2;205;203;203m█[0m[38;2;95;89;89m█[0m[38;2;246;245;245m█[0m[38;2;250;249;250m█[0m[38;2;249;247;248m█[0m[38;2;250;249;250m█[0m[38;2;238;236;236m█[0m[38;2;182;172;173m█[0m[38;2;158;145;145m█[0m[38;2;82;77;75m█[0m[38;2;140;138;141m█[0m[38;2;169;196;209m█[0m[38;2;179;225;244m█[0m[38;2;178;223;242m█[0m[38;2;177;220;239m█[0m[38;2;179;223;243m█[0m[38;2;181;229;248m█[0m[38;2;168;203;216m█[0m[38;2;77;73;77m█[0m[38;2;156;155;157m█[0m[38;2;175;175;180m█[0m[38;2;174;173;179m███[0m[38;2;176;175;181m██[0m[38;2;171;168;173m█[0m[38;2;84;78;81m█[0m[38;2;145;142;148m█[0m[38;2;181;181;187m█[0m[38;2;179;179;185m█[0m[38;2;177;175;181m█[0m[38;2;173;171;176m█[0m[38;2;169;167;172m█[0m[38;2;159;155;160m█[0m[38;2;78;73;72m█[0m[38;2;119;111;110m█[0m");
		$display("[38;2;175;174;180m█[0m[38;2;180;179;184m█[0m[38;2;110;105;108m█[0m[38;2;75;68;69m█[0m[38;2;173;172;176m█[0m[38;2;179;178;184m█[0m[38;2;179;179;184m██[0m[38;2;175;175;179m█[0m[38;2;161;154;156m█[0m[38;2;115;96;98m█[0m[38;2;69;57;58m█[0m[38;2;125;123;126m█[0m[38;2;179;180;185m█[0m[38;2;173;173;179m█[0m[38;2;174;174;179m█[0m[38;2;174;173;179m█[0m[38;2;173;172;178m█[0m[38;2;171;172;176m█[0m[38;2;175;175;178m█[0m[38;2;103;98;101m█[0m[38;2;104;99;103m█[0m[38;2;183;182;187m█[0m[38;2;178;177;183m█[0m[38;2;176;175;181m█[0m[38;2;175;174;179m█[0m[38;2;207;205;208m█[0m[38;2;225;221;221m█[0m[38;2;147;141;139m█[0m[38;2;113;107;106m█[0m[38;2;229;225;224m█[0m[38;2;234;232;233m█[0m[38;2;250;249;249m█[0m[38;2;249;248;248m█[0m[38;2;250;246;245m█[0m[38;2;255;240;242m█[0m[38;2;196;176;177m█[0m[38;2;124;108;109m█[0m[38;2;210;173;179m█[0m[38;2;100;64;68m█[0m[38;2;103;81;81m█[0m[38;2;118;103;101m█[0m[38;2;120;104;103m█[0m[38;2;115;98;96m█[0m[38;2;92;71;69m█[0m[38;2;106;85;83m█[0m[38;2;214;208;206m█[0m[38;2;255;253;254m█[0m[38;2;218;221;223m█[0m[38;2;202;224;229m█[0m[38;2;204;236;245m█[0m[38;2;205;234;243m█[0m[38;2;194;207;211m█[0m[38;2;252;251;250m█[0m[38;2;202;194;192m█[0m[38;2;98;76;77m█[0m[38;2;95;71;73m█[0m[38;2;118;99;100m█[0m[38;2;123;107;106m█[0m[38;2;121;106;103m█[0m[38;2;100;74;75m█[0m[38;2;99;66;70m█[0m[38;2;213;184;188m█[0m[38;2;210;189;191m█[0m[38;2;103;91;90m█[0m[38;2;251;231;235m█[0m[38;2;252;244;246m█[0m[38;2;250;249;248m█[0m[38;2;249;247;248m█[0m[38;2;248;246;247m█[0m[38;2;248;246;246m█[0m[38;2;234;232;229m█[0m[38;2;105;98;98m█[0m[38;2;231;226;226m█[0m[38;2;244;252;255m█[0m[38;2;189;230;245m█[0m[38;2;177;223;242m█[0m[38;2;179;224;243m█[0m[38;2;181;227;247m█[0m[38;2;180;227;246m█[0m[38;2;171;210;225m█[0m[38;2;81;80;83m█[0m[38;2;163;163;166m█[0m[38;2;180;179;185m█[0m[38;2;176;175;181m█[0m[38;2;174;173;179m██[0m[38;2;173;172;178m█[0m[38;2;175;174;180m█[0m[38;2;170;168;172m█[0m[38;2;80;74;76m█[0m[38;2;147;142;149m█[0m[38;2;180;179;185m█[0m[38;2;177;176;182m█[0m[38;2;177;176;181m█[0m[38;2;176;175;181m█[0m[38;2;173;173;179m█[0m[38;2;171;170;176m█[0m[38;2;80;75;76m█[0m[38;2;133;132;135m█[0m");
		$display("[38;2;176;175;181m█[0m[38;2;185;183;189m█[0m[38;2;112;105;108m█[0m[38;2;75;68;69m█[0m[38;2;174;172;174m█[0m[38;2;170;167;170m█[0m[38;2;155;146;151m█[0m[38;2;143;130;132m█[0m[38;2;130;110;110m█[0m[38;2;117;93;92m█[0m[38;2;148;133;133m█[0m[38;2;79;69;68m█[0m[38;2;104;92;93m█[0m[38;2;172;169;172m█[0m[38;2;175;175;180m█[0m[38;2;172;172;177m█[0m[38;2;175;174;180m█[0m[38;2;176;175;181m██[0m[38;2;180;177;182m█[0m[38;2;104;99;100m█[0m[38;2;108;104;108m█[0m[38;2;182;181;186m█[0m[38;2;178;177;182m█[0m[38;2;175;174;180m█[0m[38;2;190;189;195m█[0m[38;2;255;255;255m█[0m[38;2;243;241;241m█[0m[38;2;139;132;131m█[0m[38;2;101;95;94m█[0m[38;2;207;203;202m█[0m[38;2;247;244;245m█[0m[38;2;249;248;249m█[0m[38;2;250;244;243m█[0m[38;2;249;210;217m█[0m[38;2;218;161;171m█[0m[38;2;151;113;119m█[0m[38;2;92;73;74m█[0m[38;2;213;158;169m█[0m[38;2;212;160;169m█[0m[38;2;187;137;146m█[0m[38;2;188;141;148m█[0m[38;2;190;170;171m█[0m[38;2;198;191;191m█[0m[38;2;219;214;214m█[0m[38;2;249;247;247m█[0m[38;2;255;252;253m█[0m[38;2;242;238;239m█[0m[38;2;206;202;202m█[0m[38;2;237;237;236m█[0m[38;2;135;128;129m█[0m[38;2;185;180;181m█[0m[38;2;231;229;228m█[0m[38;2;207;202;202m█[0m[38;2;255;254;254m█[0m[38;2;248;246;246m█[0m[38;2;220;214;214m█[0m[38;2;202;194;195m█[0m[38;2;197;190;190m█[0m[38;2;204;178;182m█[0m[38;2;201;151;160m█[0m[38;2;174;125;132m█[0m[38;2;223;168;178m█[0m[38;2;156;117;124m█[0m[38;2;92;73;73m█[0m[38;2;203;150;159m█[0m[38;2;226;175;183m█[0m[38;2;239;211;215m█[0m[38;2;250;248;248m█[0m[38;2;251;250;251m█[0m[38;2;218;214;214m█[0m[38;2;169;161;160m█[0m[38;2;92;82;82m█[0m[38;2;133;121;122m█[0m[38;2;165;152;151m█[0m[38;2;169;188;196m█[0m[38;2;177;223;241m█[0m[38;2;175;217;234m█[0m[38;2;135;156;167m█[0m[38;2;117;125;135m█[0m[38;2;114;119;127m█[0m[38;2;75;69;72m█[0m[38;2;146;142;145m█[0m[38;2;181;180;186m█[0m[38;2;179;178;184m█[0m[38;2;176;175;181m█[0m[38;2;173;173;178m██[0m[38;2;177;176;182m█[0m[38;2;174;171;177m█[0m[38;2;84;78;82m█[0m[38;2;145;141;146m█[0m[38;2;178;177;183m█[0m[38;2;179;178;183m█[0m[38;2;166;163;168m█[0m[38;2;158;151;155m█[0m[38;2;158;154;160m█[0m[38;2;172;171;177m█[0m[38;2;83;77;78m█[0m[38;2;127;125;128m█[0m");
		$display("[38;2;174;170;176m█[0m[38;2;169;161;165m█[0m[38;2;104;95;96m█[0m[38;2;70;61;60m█[0m[38;2;134;120;119m█[0m[38;2;141;128;129m█[0m[38;2;151;141;144m█[0m[38;2;168;164;166m█[0m[38;2;167;161;163m█[0m[38;2;146;135;137m█[0m[38;2;158;147;150m█[0m[38;2;79;70;69m█[0m[38;2;111;101;102m█[0m[38;2;124;105;107m█[0m[38;2;164;159;161m█[0m[38;2;178;178;184m█[0m[38;2;177;176;182m█[0m[38;2;179;178;184m█[0m[38;2;181;180;186m█[0m[38;2;182;178;183m█[0m[38;2;102;97;100m█[0m[38;2;115;113;114m█[0m[38;2;182;181;186m█[0m[38;2;176;175;181m█[0m[38;2;173;173;179m█[0m[38;2;188;186;190m█[0m[38;2;169;158;160m█[0m[38;2;162;149;149m█[0m[38;2;130;121;121m█[0m[38;2;119;115;113m█[0m[38;2;234;232;232m█[0m[38;2;248;245;246m█[0m[38;2;249;249;249m█[0m[38;2;249;240;240m█[0m[38;2;248;194;203m█[0m[38;2;211;154;162m█[0m[38;2;182;143;147m█[0m[38;2;104;83;83m█[0m[38;2;220;164;172m█[0m[38;2;231;173;182m█[0m[38;2;226;168;177m█[0m[38;2;252;196;205m█[0m[38;2;255;239;242m█[0m[38;2;255;255;255m█[0m[38;2;253;251;252m█[0m[38;2;250;248;249m█[0m[38;2;249;248;249m█[0m[38;2;247;245;246m█[0m[38;2;189;183;183m█[0m[38;2;171;162;162m█[0m[38;2;162;150;149m█[0m[38;2;155;144;142m█[0m[38;2;173;162;161m█[0m[38;2;212;206;205m█[0m[38;2;251;250;249m█[0m[38;2;250;248;249m█[0m[38;2;253;251;252m█[0m[38;2;254;253;254m█[0m[38;2;255;255;255m█[0m[38;2;255;219;230m█[0m[38;2;228;167;178m█[0m[38;2;234;175;183m█[0m[38;2;225;167;177m█[0m[38;2;168;129;136m█[0m[38;2;93;72;73m█[0m[38;2;222;167;174m█[0m[38;2;210;152;161m█[0m[38;2;241;201;208m█[0m[38;2;250;247;247m█[0m[38;2;249;247;249m█[0m[38;2;251;250;251m█[0m[38;2;255;254;255m█[0m[38;2;112;105;107m█[0m[38;2;205;202;201m█[0m[38;2;224;219;217m█[0m[38;2;165;179;187m█[0m[38;2;173;217;235m█[0m[38;2;177;221;239m█[0m[38;2;168;208;225m█[0m[38;2;175;216;234m█[0m[38;2;155;188;201m█[0m[38;2;73;67;71m█[0m[38;2;146;141;144m█[0m[38;2;181;180;186m█[0m[38;2;180;180;185m██[0m[38;2;178;177;183m█[0m[38;2;176;175;181m█[0m[38;2;178;178;184m█[0m[38;2;179;176;181m█[0m[38;2;89;84;87m█[0m[38;2;143;140;142m█[0m[38;2;180;179;185m█[0m[38;2;179;179;184m█[0m[38;2;180;178;183m█[0m[38;2;175;173;178m█[0m[38;2;178;176;182m█[0m[38;2;173;173;178m█[0m[38;2;83;78;78m█[0m[38;2;116;114;115m█[0m");
		$display("[38;2;134;116;117m█[0m[38;2;144;127;128m█[0m[38;2;106;98;97m█[0m[38;2;72;67;67m█[0m[38;2;171;167;171m█[0m[38;2;181;181;187m█[0m[38;2;183;184;189m█[0m[38;2;184;184;190m█[0m[38;2;184;183;189m█[0m[38;2;174;170;175m█[0m[38;2;164;158;161m█[0m[38;2;88;82;83m█[0m[38;2;128;127;129m█[0m[38;2;167;161;163m█[0m[38;2;118;98;99m█[0m[38;2;161;153;157m█[0m[38;2;182;182;188m██[0m[38;2;182;181;187m█[0m[38;2;183;181;185m█[0m[38;2;99;95;95m█[0m[38;2;125;124;125m█[0m[38;2;184;184;188m█[0m[38;2;178;178;183m█[0m[38;2;179;179;185m█[0m[38;2;167;164;168m█[0m[38;2;191;183;185m█[0m[38;2;255;255;255m█[0m[38;2;176;174;172m█[0m[38;2;123;118;118m█[0m[38;2;230;227;227m█[0m[38;2;242;239;240m█[0m[38;2;250;248;249m█[0m[38;2;249;247;248m█[0m[38;2;249;235;237m█[0m[38;2;255;225;228m█[0m[38;2;192;162;166m█[0m[38;2;90;75;74m█[0m[38;2;245;202;209m█[0m[38;2;254;213;219m█[0m[38;2;253;221;226m█[0m[38;2;249;236;236m█[0m[38;2;249;248;246m█[0m[38;2;249;247;248m█████[0m[38;2;255;255;255m█[0m[38;2;242;239;240m█[0m[38;2;209;202;202m█[0m[38;2;203;198;197m█[0m[38;2;238;237;237m█[0m[38;2;254;254;253m█[0m[38;2;249;247;248m████[0m[38;2;250;247;248m█[0m[38;2;250;244;246m█[0m[38;2;252;226;232m█[0m[38;2;253;212;218m█[0m[38;2;255;210;219m█[0m[38;2;196;162;167m█[0m[38;2;119;99;101m█[0m[38;2;255;214;221m█[0m[38;2;253;223;228m█[0m[38;2;249;241;243m█[0m[38;2;249;248;248m█[0m[38;2;251;249;250m█[0m[38;2;234;231;232m█[0m[38;2;178;169;171m█[0m[38;2;93;84;85m█[0m[38;2;170;162;159m█[0m[38;2;247;248;247m█[0m[38;2;196;234;249m█[0m[38;2;177;223;243m█[0m[38;2;177;221;241m█[0m[38;2;172;213;231m█[0m[38;2;174;216;234m█[0m[38;2;158;191;205m█[0m[38;2;80;74;77m█[0m[38;2;174;174;176m█[0m[38;2;181;180;186m█[0m[38;2;179;179;185m█[0m[38;2;181;180;186m██[0m[38;2;180;179;185m█[0m[38;2;181;181;186m█[0m[38;2;186;184;187m█[0m[38;2;97;93;96m█[0m[38;2;136;132;135m█[0m[38;2;188;186;191m█[0m[38;2;182;181;187m█[0m[38;2;181;180;186m█[0m[38;2;182;181;187m█[0m[38;2;180;180;185m█[0m[38;2;176;176;181m█[0m[38;2;79;76;75m█[0m[38;2;108;105;107m█[0m");
		$display("[38;2;182;181;187m█[0m[38;2;189;187;192m█[0m[38;2;130;126;128m█[0m[38;2;69;65;66m█[0m[38;2;173;170;175m█[0m[38;2;180;180;185m██[0m[38;2;182;181;187m█[0m[38;2;181;180;186m█[0m[38;2;182;181;186m█[0m[38;2;184;184;187m█[0m[38;2;93;88;92m█[0m[38;2;123;117;123m█[0m[38;2;186;186;191m█[0m[38;2;169;163;166m█[0m[38;2;132;115;116m█[0m[38;2;146;133;136m█[0m[38;2;174;168;172m█[0m[38;2;184;183;188m█[0m[38;2;190;189;193m█[0m[38;2;100;96;97m█[0m[38;2;134;132;135m█[0m[38;2;189;189;194m█[0m[38;2;182;182;188m█[0m[38;2;181;182;187m█[0m[38;2;181;181;187m█[0m[38;2;212;211;216m█[0m[38;2;246;244;244m█[0m[38;2;138;129;129m█[0m[38;2;94;85;85m█[0m[38;2;193;187;185m█[0m[38;2;241;239;240m█[0m[38;2;255;253;254m█[0m[38;2;249;247;248m█[0m[38;2;251;251;251m█[0m[38;2;255;254;255m█[0m[38;2;205;200;201m█[0m[38;2;78;74;73m█[0m[38;2;234;232;231m█[0m[38;2;251;251;251m█[0m[38;2;250;249;250m█[0m[38;2;249;249;249m█[0m[38;2;249;247;248m███████[0m[38;2;250;248;249m█[0m[38;2;253;252;253m██[0m[38;2;250;248;249m█[0m[38;2;249;247;248m██████[0m[38;2;249;248;249m█[0m[38;2;249;249;250m█[0m[38;2;249;249;249m█[0m[38;2;255;253;254m█[0m[38;2;189;185;186m█[0m[38;2;124;117;118m█[0m[38;2;255;252;252m█[0m[38;2;248;249;248m█[0m[38;2;251;250;251m█[0m[38;2;253;252;253m█[0m[38;2;249;247;248m█[0m[38;2;247;245;246m█[0m[38;2;246;244;245m█[0m[38;2;130;122;124m█[0m[38;2;120;111;110m█[0m[38;2;136;138;144m█[0m[38;2;169;206;224m█[0m[38;2;181;227;248m█[0m[38;2;167;206;222m█[0m[38;2;133;151;161m█[0m[38;2;126;136;146m█[0m[38;2;112;114;120m█[0m[38;2;81;75;77m█[0m[38;2;170;170;173m█[0m[38;2;183;182;188m█[0m[38;2;182;181;187m██[0m[38;2;184;183;189m██[0m[38;2;183;182;188m█[0m[38;2;188;188;191m█[0m[38;2;108;104;106m█[0m[38;2;128;124;126m█[0m[38;2;190;188;192m█[0m[38;2;182;181;187m█[0m[38;2;179;178;184m█[0m[38;2;179;179;185m█[0m[38;2;182;181;187m█[0m[38;2;178;177;182m█[0m[38;2;79;75;75m█[0m[38;2;109;106;109m█[0m");
		$display("[38;2;185;184;190m█[0m[38;2;188;186;191m█[0m[38;2;133;131;132m█[0m[38;2;67;63;64m█[0m[38;2;173;170;176m█[0m[38;2;183;184;189m█[0m[38;2;180;179;185m██[0m[38;2;182;181;187m█[0m[38;2;183;182;187m█[0m[38;2;185;184;187m█[0m[38;2;96;88;91m█[0m[38;2;117;114;116m█[0m[38;2;188;188;192m█[0m[38;2;185;185;190m█[0m[38;2;186;184;188m█[0m[38;2;161;150;152m█[0m[38;2;137;121;121m█[0m[38;2;136;119;121m█[0m[38;2;146;130;132m█[0m[38;2;92;81;83m█[0m[38;2;122;116;117m█[0m[38;2;166;159;163m█[0m[38;2;168;162;166m█[0m[38;2;173;170;174m█[0m[38;2;178;174;179m█[0m[38;2;186;183;188m█[0m[38;2;166;157;159m█[0m[38;2;78;65;66m█[0m[38;2;134;130;129m█[0m[38;2;255;255;255m█[0m[38;2;232;228;229m█[0m[38;2;212;207;208m█[0m[38;2;255;254;254m█[0m[38;2;237;233;234m█[0m[38;2;254;251;251m█[0m[38;2;229;226;224m█[0m[38;2;79;75;74m█[0m[38;2;227;225;224m█[0m[38;2;255;255;255m█[0m[38;2;252;249;250m█[0m[38;2;250;247;248m█[0m[38;2;249;247;248m████████████████████[0m[38;2;255;255;255m█[0m[38;2;182;179;180m█[0m[38;2;123;120;118m█[0m[38;2;255;255;255m█[0m[38;2;255;254;255m█[0m[38;2;239;237;237m█[0m[38;2;213;209;210m█[0m[38;2;244;241;241m█[0m[38;2;177;168;168m█[0m[38;2;200;193;194m█[0m[38;2;153;148;150m█[0m[38;2;133;150;159m█[0m[38;2;182;224;242m█[0m[38;2;176;219;238m█[0m[38;2;181;228;247m█[0m[38;2;182;229;249m█[0m[38;2;182;230;249m█[0m[38;2;183;230;249m█[0m[38;2;159;178;185m█[0m[38;2;74;70;71m█[0m[38;2;166;164;167m█[0m[38;2;184;183;189m█[0m[38;2;182;181;187m█[0m[38;2;182;181;188m█[0m[38;2;180;179;185m█[0m[38;2;183;182;188m█[0m[38;2;184;183;189m█[0m[38;2;191;188;193m█[0m[38;2;115;110;114m██[0m[38;2;186;186;190m█[0m[38;2;180;180;186m█[0m[38;2;181;180;186m█[0m[38;2;180;181;186m█[0m[38;2;183;182;188m█[0m[38;2;181;179;185m█[0m[38;2;82;77;77m█[0m[38;2;119;116;116m█[0m");
		$display("[38;2;184;183;189m█[0m[38;2;190;188;194m█[0m[38;2;140;137;140m█[0m[38;2;67;62;64m█[0m[38;2;172;170;174m█[0m[38;2;186;186;191m█[0m[38;2;185;184;190m█[0m[38;2;184;183;189m█[0m[38;2;182;181;187m█[0m[38;2;181;181;186m█[0m[38;2;182;181;185m█[0m[38;2;92;84;88m█[0m[38;2;121;119;121m█[0m[38;2;189;189;194m█[0m[38;2;185;184;189m█[0m[38;2;185;184;190m█[0m[38;2;188;187;193m█[0m[38;2;188;187;192m█[0m[38;2;182;180;184m█[0m[38;2;176;170;174m█[0m[38;2;92;85;85m█[0m[38;2;119;110;111m█[0m[38;2;156;144;145m█[0m[38;2;135;118;116m█[0m[38;2;106;80;78m█[0m[38;2;130;106;106m█[0m[38;2;132;113;114m█[0m[38;2;141;126;126m█[0m[38;2;104;93;93m█[0m[38;2;127;121;121m█[0m[38;2;228;226;225m█[0m[38;2;134;122;124m█[0m[38;2;217;211;212m█[0m[38;2;188;178;177m█[0m[38;2;94;73;71m█[0m[38;2;149;132;130m█[0m[38;2;161;149;147m█[0m[38;2;101;93;89m█[0m[38;2;167;157;156m█[0m[38;2;179;170;170m█[0m[38;2;236;232;231m█[0m[38;2;255;253;252m█[0m[38;2;255;253;254m█[0m[38;2;255;254;255m█[0m[38;2;255;253;254m█[0m[38;2;254;252;253m█[0m[38;2;253;252;253m█[0m[38;2;252;251;252m█[0m[38;2;252;250;251m██[0m[38;2;251;250;251m██[0m[38;2;252;250;251m██[0m[38;2;252;251;252m█[0m[38;2;253;251;253m█[0m[38;2;254;252;254m█[0m[38;2;255;253;255m█[0m[38;2;255;254;255m██[0m[38;2;253;252;253m█[0m[38;2;252;250;250m█[0m[38;2;171;162;162m█[0m[38;2;165;154;153m█[0m[38;2;140;131;129m█[0m[38;2;177;168;167m█[0m[38;2;156;142;142m█[0m[38;2;101;80;79m█[0m[38;2;87;67;66m█[0m[38;2;204;216;221m█[0m[38;2;200;227;238m█[0m[38;2;132;146;152m█[0m[38;2;97;92;95m█[0m[38;2;114;132;144m█[0m[38;2;184;231;251m█[0m[38;2;175;218;236m█[0m[38;2;147;172;188m█[0m[38;2;143;166;180m█[0m[38;2;161;197;212m█[0m[38;2;184;219;234m█[0m[38;2;166;169;172m█[0m[38;2;81;75;76m█[0m[38;2;174;172;177m█[0m[38;2;186;185;191m█[0m[38;2;183;181;186m█[0m[38;2;160;155;159m█[0m[38;2;181;180;185m█[0m[38;2;183;182;188m█[0m[38;2;184;184;189m█[0m[38;2;189;186;191m█[0m[38;2;116;112;114m█[0m[38;2;106;102;104m█[0m[38;2;188;187;192m█[0m[38;2;183;182;188m█[0m[38;2;185;184;189m█[0m[38;2;183;182;188m█[0m[38;2;184;183;189m█[0m[38;2;183;183;188m█[0m[38;2;89;83;85m█[0m[38;2;89;73;72m█[0m");
		$display("[38;2;186;186;191m█[0m[38;2;191;191;196m█[0m[38;2;138;134;138m█[0m[38;2;70;65;67m█[0m[38;2;177;175;180m█[0m[38;2;187;186;192m█[0m[38;2;188;187;192m█[0m[38;2;188;187;193m█[0m[38;2;186;185;191m█[0m[38;2;185;185;190m█[0m[38;2;181;181;184m█[0m[38;2;82;77;80m█[0m[38;2;135;130;133m█[0m[38;2;190;189;194m█[0m[38;2;186;185;190m█[0m[38;2;186;185;191m█[0m[38;2;189;188;193m█[0m[38;2;189;188;194m█[0m[38;2;188;187;193m█[0m[38;2;191;189;195m█[0m[38;2;95;88;89m█[0m[38;2;137;134;137m█[0m[38;2;195;198;202m█[0m[38;2;185;184;188m█[0m[38;2;119;98;98m█[0m[38;2;164;154;155m█[0m[38;2;183;181;186m█[0m[38;2;184;182;188m█[0m[38;2;113;110;111m█[0m[38;2;106;102;101m█[0m[38;2;180;177;180m█[0m[38;2;175;173;177m█[0m[38;2;197;195;199m█[0m[38;2;66;42;42m█[0m[38;2;160;145;141m█[0m[38;2;121;101;98m█[0m[38;2;105;83;83m█[0m[38;2;245;242;240m█[0m[38;2;255;254;253m█[0m[38;2;157;146;145m█[0m[38;2;185;175;174m█[0m[38;2;198;191;190m█[0m[38;2;181;170;170m█[0m[38;2;190;180;180m█[0m[38;2;197;189;189m█[0m[38;2;206;198;198m█[0m[38;2;213;207;206m█[0m[38;2;219;213;212m█[0m[38;2;224;218;217m█[0m[38;2;227;221;220m█[0m[38;2;230;225;224m█[0m[38;2;231;226;226m█[0m[38;2;226;222;221m█[0m[38;2;223;219;219m█[0m[38;2;219;214;214m█[0m[38;2;212;206;206m█[0m[38;2;204;197;197m█[0m[38;2;197;189;189m█[0m[38;2;183;173;174m█[0m[38;2;173;161;162m█[0m[38;2;178;166;168m█[0m[38;2;197;187;187m█[0m[38;2;134;120;120m█[0m[38;2;247;247;243m█[0m[38;2;255;255;255m█[0m[38;2;124;108;106m█[0m[38;2;108;85;84m█[0m[38;2;166;150;147m█[0m[38;2;50;18;15m█[0m[38;2;140;161;173m█[0m[38;2;180;230;250m█[0m[38;2;184;233;251m█[0m[38;2;124;143;151m█[0m[38;2;104;119;129m█[0m[38;2;185;232;251m█[0m[38;2;181;227;245m█[0m[38;2;166;202;217m█[0m[38;2;148;176;190m█[0m[38;2;122;128;136m█[0m[38;2;121;113;115m█[0m[38;2;164;160;163m█[0m[38;2;84;80;82m█[0m[38;2;176;174;178m█[0m[38;2;189;188;193m█[0m[38;2;178;175;179m█[0m[38;2;169;161;164m█[0m[38;2;160;150;154m█[0m[38;2;178;173;178m█[0m[38;2;173;168;173m█[0m[38;2;188;187;192m█[0m[38;2;112;109;110m█[0m[38;2;103;101;101m█[0m[38;2;188;187;193m█[0m[38;2;185;184;190m█[0m[38;2;186;185;191m█[0m[38;2;186;185;190m█[0m[38;2;188;188;193m█[0m[38;2;176;173;176m█[0m[38;2;86;77;78m█[0m[38;2;109;102;102m█[0m");
		$display("[38;2;188;187;193m█[0m[38;2;193;192;199m█[0m[38;2;136;132;136m█[0m[38;2;77;71;73m█[0m[38;2;170;165;168m█[0m[38;2;167;162;166m█[0m[38;2;190;188;194m█[0m[38;2;164;157;164m█[0m[38;2;186;183;189m█[0m[38;2;188;187;193m█[0m[38;2;179;179;183m█[0m[38;2;77;72;75m█[0m[38;2;147;141;145m█[0m[38;2;192;191;196m█[0m[38;2;189;188;194m█[0m[38;2;190;189;195m█[0m[38;2;191;190;196m██[0m[38;2;190;189;195m█[0m[38;2;191;190;195m█[0m[38;2;94;88;88m█[0m[38;2;140;136;140m█[0m[38;2;191;192;197m█[0m[38;2;190;191;195m█[0m[38;2;154;141;141m█[0m[38;2;130;109;109m█[0m[38;2;190;189;193m█[0m[38;2;192;191;197m█[0m[38;2;125;121;122m█[0m[38;2;105;100;101m█[0m[38;2;191;190;194m█[0m[38;2;190;189;196m█[0m[38;2;187;186;192m█[0m[38;2;131;119;120m█[0m[38;2;114;95;92m█[0m[38;2;83;57;54m█[0m[38;2;86;61;59m█[0m[38;2;202;196;191m█[0m[38;2;213;207;204m█[0m[38;2;96;75;75m█[0m[38;2;133;115;114m█[0m[38;2;179;167;164m█[0m[38;2;180;167;165m█[0m[38;2;136;124;122m█[0m[38;2;162;149;148m█[0m[38;2;170;155;154m█[0m[38;2;166;151;149m█[0m[38;2;162;147;145m█[0m[38;2;159;143;141m█[0m[38;2;156;141;137m█[0m[38;2;142;127;122m█[0m[38;2;128;113;110m█[0m[38;2;146;133;129m█[0m[38;2;147;131;129m█[0m[38;2;148;133;131m█[0m[38;2;152;138;136m█[0m[38;2;162;147;146m█[0m[38;2;127;113;113m█[0m[38;2;175;163;162m█[0m[38;2;192;183;181m█[0m[38;2;196;186;185m█[0m[38;2;164;149;148m█[0m[38;2;97;73;74m█[0m[38;2;204;195;193m█[0m[38;2;202;194;193m█[0m[38;2;91;67;66m█[0m[38;2;92;66;62m█[0m[38;2;106;88;85m█[0m[38;2;114;119;126m█[0m[38;2;177;217;236m█[0m[38;2;179;225;244m█[0m[38;2;184;232;250m█[0m[38;2;129;152;160m█[0m[38;2;95;104;110m█[0m[38;2;146;169;182m█[0m[38;2;137;157;167m█[0m[38;2;166;202;219m█[0m[38;2;188;227;244m█[0m[38;2;187;199;206m█[0m[38;2;172;166;170m█[0m[38;2;165;158;162m█[0m[38;2;84;79;83m█[0m[38;2;177;175;178m█[0m[38;2;186;185;190m█[0m[38;2;185;186;190m█[0m[38;2;188;189;193m█[0m[38;2;176;171;177m█[0m[38;2;185;180;186m█[0m[38;2;177;170;177m█[0m[38;2;196;193;199m█[0m[38;2;110;105;107m█[0m[38;2;111;108;108m█[0m[38;2;191;188;195m█[0m[38;2;183;182;188m█[0m[38;2;186;186;192m█[0m[38;2;189;189;194m█[0m[38;2;161;152;155m█[0m[38;2;121;100;100m█[0m[38;2;77;67;65m█[0m[38;2;129;128;129m█[0m");
		$display("[38;2;188;187;193m█[0m[38;2;194;193;199m█[0m[38;2;132;129;132m█[0m[38;2;81;76;78m█[0m[38;2;176;173;175m█[0m[38;2;157;149;151m█[0m[38;2;177;171;176m█[0m[38;2;174;170;177m█[0m[38;2;184;183;189m█[0m[38;2;186;185;191m█[0m[38;2;180;180;183m█[0m[38;2;76;70;73m█[0m[38;2;137;134;136m█[0m[38;2;188;188;193m█[0m[38;2;186;185;190m█[0m[38;2;190;189;195m██[0m[38;2;188;187;193m█[0m[38;2;189;188;195m█[0m[38;2;191;191;196m█[0m[38;2;93;86;88m█[0m[38;2;136;131;136m█[0m[38;2;189;188;194m█[0m[38;2;187;188;193m█[0m[38;2;169;154;155m█[0m[38;2;124;101;99m█[0m[38;2;193;193;198m█[0m[38;2;195;194;200m█[0m[38;2;134;131;134m█[0m[38;2;101;98;98m█[0m[38;2;191;190;193m█[0m[38;2;190;189;194m█[0m[38;2;189;188;194m█[0m[38;2;190;189;194m█[0m[38;2;177;170;175m█[0m[38;2;93;70;70m█[0m[38;2;80;55;54m█[0m[38;2;87;73;70m█[0m[38;2;91;74;69m█[0m[38;2;82;57;54m█[0m[38;2;76;48;46m█[0m[38;2;69;40;39m█[0m[38;2;72;44;43m█[0m[38;2;73;59;56m█[0m[38;2;76;56;54m█[0m[38;2;85;59;55m█[0m[38;2;89;63;60m█[0m[38;2;93;68;66m█[0m[38;2;97;73;71m█[0m[38;2;100;75;74m█[0m[38;2;98;81;78m█[0m[38;2;87;76;73m█[0m[38;2;107;86;85m█[0m[38;2;106;81;79m█[0m[38;2;101;78;74m█[0m[38;2;98;76;73m█[0m[38;2;99;77;76m█[0m[38;2;82;69;67m█[0m[38;2;79;59;57m█[0m[38;2;73;46;44m█[0m[38;2;64;35;35m█[0m[38;2;63;33;33m█[0m[38;2;69;40;41m█[0m[38;2;83;62;61m█[0m[38;2;81;64;63m█[0m[38;2;130;111;109m█[0m[38;2;89;63;59m█[0m[38;2;105;104;109m█[0m[38;2;187;235;255m█[0m[38;2;179;225;246m█[0m[38;2;174;217;236m█[0m[38;2;176;217;234m█[0m[38;2;130;150;159m█[0m[38;2;101;113;118m█[0m[38;2;180;222;243m█[0m[38;2;158;184;195m█[0m[38;2;112;107;114m█[0m[38;2;152;148;152m█[0m[38;2;191;189;193m█[0m[38;2;198;197;203m█[0m[38;2;174;171;175m█[0m[38;2;84;80;81m█[0m[38;2;182;181;186m█[0m[38;2;188;188;194m█[0m[38;2;186;185;191m█[0m[38;2;187;186;191m█[0m[38;2;189;188;193m█[0m[38;2;190;189;195m█[0m[38;2;192;191;197m█[0m[38;2;196;193;199m█[0m[38;2;106;101;103m█[0m[38;2;126;123;123m█[0m[38;2;193;193;199m█[0m[38;2;190;191;196m█[0m[38;2;179;173;177m█[0m[38;2;137;118;120m█[0m[38;2;131;108;110m█[0m[38;2;176;167;168m█[0m[38;2;86;83;83m█[0m[38;2;127;125;127m█[0m");
		$display("[38;2;186;185;190m█[0m[38;2;191;191;196m█[0m[38;2;125;120;122m█[0m[38;2;88;83;84m█[0m[38;2;192;193;195m█[0m[38;2;180;176;180m█[0m[38;2;190;188;193m█[0m[38;2;191;191;197m█[0m[38;2;191;190;196m█[0m[38;2;192;191;197m█[0m[38;2;186;184;188m█[0m[38;2;79;72;75m█[0m[38;2;134;132;135m█[0m[38;2;193;194;198m█[0m[38;2;189;188;194m█[0m[38;2;191;190;196m█[0m[38;2;192;191;197m█[0m[38;2;191;190;196m██[0m[38;2;195;194;198m█[0m[38;2;96;89;91m█[0m[38;2;128;122;127m█[0m[38;2;193;191;197m█[0m[38;2;192;193;198m█[0m[38;2;153;140;141m█[0m[38;2;137;119;118m█[0m[38;2;198;197;203m█[0m[38;2;194;191;196m█[0m[38;2;117;108;111m█[0m[38;2;100;97;98m█[0m[38;2;192;189;192m█[0m[38;2;188;187;192m█[0m[38;2;188;187;193m██[0m[38;2;192;193;199m█[0m[38;2;159;149;152m█[0m[38;2;77;53;52m█[0m[38;2;82;69;66m█[0m[38;2;172;165;164m█[0m[38;2;241;236;235m█[0m[38;2;239;233;232m█[0m[38;2;234;228;228m█[0m[38;2;230;223;223m█[0m[38;2;106;98;97m█[0m[38;2;167;158;157m█[0m[38;2;207;197;196m█[0m[38;2;190;177;175m█[0m[38;2;182;168;167m█[0m[38;2;173;159;157m█[0m[38;2;167;155;154m█[0m[38;2;132;122;120m█[0m[38;2;93;82;82m█[0m[38;2;179;164;164m█[0m[38;2;175;161;159m█[0m[38;2;168;154;152m█[0m[38;2;166;152;151m█[0m[38;2;162;151;147m█[0m[38;2;80;72;70m█[0m[38;2;164;152;152m█[0m[38;2;199;188;186m█[0m[38;2;209;199;197m█[0m[38;2;219;212;211m█[0m[38;2;232;226;226m█[0m[38;2;198;194;194m█[0m[38;2;119;113;112m█[0m[38;2;203;193;190m█[0m[38;2;87;68;68m█[0m[38;2;158;185;200m█[0m[38;2;179;227;244m█[0m[38;2;181;228;245m█[0m[38;2;171;212;230m█[0m[38;2;127;141;149m█[0m[38;2;87;84;86m█[0m[38;2;112;120;126m█[0m[38;2;189;217;230m█[0m[38;2;193;201;210m█[0m[38;2;189;188;192m█[0m[38;2;166;156;158m█[0m[38;2;151;135;138m█[0m[38;2;155;139;141m█[0m[38;2;140;127;129m█[0m[38;2;82;75;75m█[0m[38;2;171;166;170m█[0m[38;2;191;187;193m█[0m[38;2;192;191;196m█[0m[38;2;189;189;194m█[0m[38;2;188;188;193m█[0m[38;2;186;185;190m█[0m[38;2;185;185;190m█[0m[38;2;193;190;195m█[0m[38;2;104;99;101m█[0m[38;2;139;137;137m█[0m[38;2;182;177;181m█[0m[38;2;144;127;130m█[0m[38;2;128;107;104m█[0m[38;2;162;149;150m█[0m[38;2;192;190;194m█[0m[38;2;188;187;189m█[0m[38;2;83;81;81m█[0m[38;2;126;124;127m█[0m");
		$display("[38;2;190;189;195m█[0m[38;2;194;195;200m█[0m[38;2;118;114;115m█[0m[38;2;96;91;91m█[0m[38;2;195;196;199m█[0m[38;2;193;192;197m█[0m[38;2;191;190;196m█[0m[38;2;192;191;197m██[0m[38;2;194;194;199m█[0m[38;2;192;188;193m█[0m[38;2;82;75;78m█[0m[38;2;145;143;145m█[0m[38;2;198;198;203m█[0m[38;2;194;192;198m█[0m[38;2;191;189;195m█[0m[38;2;179;176;180m█[0m[38;2;170;164;167m█[0m[38;2;190;188;192m█[0m[38;2;197;197;202m█[0m[38;2;103;97;99m█[0m[38;2;133;128;132m█[0m[38;2;200;198;204m█[0m[38;2;198;197;202m█[0m[38;2;134;113;117m█[0m[38;2;157;143;144m█[0m[38;2;194;195;200m█[0m[38;2;188;186;191m█[0m[38;2;124;114;116m█[0m[38;2;97;90;91m█[0m[38;2;178;174;178m█[0m[38;2;191;189;195m█[0m[38;2;192;191;197m██[0m[38;2;192;191;196m█[0m[38;2;196;195;200m█[0m[38;2;130;118;120m█[0m[38;2;68;56;54m█[0m[38;2;77;57;57m█[0m[38;2;104;81;81m█[0m[38;2;121;99;102m█[0m[38;2;136;117;116m█[0m[38;2;146;129;126m█[0m[38;2;92;80;79m█[0m[38;2;132;120;118m█[0m[38;2;180;167;166m█[0m[38;2;200;188;188m█[0m[38;2;209;199;198m█[0m[38;2;213;203;202m█[0m[38;2;218;210;209m█[0m[38;2;165;158;157m█[0m[38;2;100;92;91m█[0m[38;2;211;201;201m█[0m[38;2;208;199;198m█[0m[38;2;207;198;197m█[0m[38;2;208;198;196m█[0m[38;2;196;188;185m█[0m[38;2;85;76;76m█[0m[38;2;160;149;148m█[0m[38;2;188;174;173m█[0m[38;2;177;162;160m█[0m[38;2;160;145;143m█[0m[38;2;135;118;115m█[0m[38;2;107;90;88m█[0m[38;2;70;55;54m█[0m[38;2;62;38;37m█[0m[38;2;124;131;137m█[0m[38;2;183;230;249m█[0m[38;2;158;191;205m█[0m[38;2;123;134;144m█[0m[38;2;184;224;240m█[0m[38;2;185;217;231m█[0m[38;2;111;109;114m█[0m[38;2;108;104;106m█[0m[38;2;198;197;201m█[0m[38;2;193;191;196m█[0m[38;2;192;191;196m█[0m[38;2;191;190;194m█[0m[38;2;189;188;192m█[0m[38;2;191;188;192m█[0m[38;2;164;159;161m█[0m[38;2;86;76;77m█[0m[38;2;153;139;141m█[0m[38;2;146;129;130m█[0m[38;2;146;128;129m█[0m[38;2;167;159;164m█[0m[38;2;188;185;190m█[0m[38;2;191;191;196m█[0m[38;2;189;188;194m█[0m[38;2;182;180;184m█[0m[38;2;101;91;93m█[0m[38;2;108;91;92m█[0m[38;2;142;120;120m█[0m[38;2;162;151;153m█[0m[38;2;189;188;191m█[0m[38;2;194;194;199m█[0m[38;2;191;192;197m█[0m[38;2;189;187;190m█[0m[38;2;84;79;79m█[0m[38;2;131;128;129m█[0m");
		$display("[38;2;193;192;198m█[0m[38;2;197;196;202m█[0m[38;2;111;105;108m█[0m[38;2;101;98;99m█[0m[38;2;196;197;199m█[0m[38;2;192;191;196m█[0m[38;2;192;191;197m██[0m[38;2;193;192;198m█[0m[38;2;195;194;200m█[0m[38;2;190;188;193m█[0m[38;2;85;78;79m█[0m[38;2;162;160;161m█[0m[38;2;200;200;205m█[0m[38;2;196;195;201m█[0m[38;2;194;193;198m█[0m[38;2;166;159;163m█[0m[38;2;182;178;182m█[0m[38;2;191;189;194m█[0m[38;2;199;199;203m█[0m[38;2;111;105;108m█[0m[38;2;140;134;139m█[0m[38;2;202;201;206m█[0m[38;2;197;194;199m█[0m[38;2;125;98;100m█[0m[38;2;174;163;164m█[0m[38;2;194;195;200m█[0m[38;2;196;195;201m█[0m[38;2;143;139;142m█[0m[38;2;88;79;82m█[0m[38;2;197;195;201m█[0m[38;2;195;194;200m█[0m[38;2;193;192;198m█[0m[38;2;194;193;198m█[0m[38;2;195;194;199m█[0m[38;2;194;193;199m█[0m[38;2;197;195;200m█[0m[38;2;104;97;99m█[0m[38;2;63;42;41m█[0m[38;2;112;91;88m█[0m[38;2;147;130;130m█[0m[38;2;131;110;108m█[0m[38;2;112;92;88m█[0m[38;2;81;70;67m█[0m[38;2;67;49;47m█[0m[38;2;67;39;36m█[0m[38;2;66;36;34m█[0m[38;2;66;37;35m█[0m[38;2;67;38;35m█[0m[38;2;66;36;38m█[0m[38;2;70;48;48m█[0m[38;2;68;55;51m█[0m[38;2;61;34;33m█[0m[38;2;63;35;32m█[0m[38;2;65;37;35m█[0m[38;2;68;40;38m█[0m[38;2;75;50;47m█[0m[38;2;73;60;57m█[0m[38;2;73;54;50m█[0m[38;2;85;61;58m█[0m[38;2;94;69;66m█[0m[38;2;103;80;76m█[0m[38;2;93;69;65m█[0m[38;2;65;40;37m█[0m[38;2;79;68;68m█[0m[38;2;140;151;157m█[0m[38;2;97;93;97m█[0m[38;2;177;200;212m█[0m[38;2;172;190;198m█[0m[38;2;84;68;69m█[0m[38;2;187;187;195m█[0m[38;2;196;196;203m█[0m[38;2;112;106;107m█[0m[38;2;122;117;119m█[0m[38;2;201;200;204m█[0m[38;2;192;191;197m█[0m[38;2;190;189;195m█[0m[38;2;189;188;194m█[0m[38;2;193;193;198m█[0m[38;2;200;199;205m█[0m[38;2;175;175;177m█[0m[38;2;90;85;86m█[0m[38;2;190;191;194m█[0m[38;2;192;191;196m█[0m[38;2;178;168;173m█[0m[38;2;150;135;137m█[0m[38;2;141;123;125m█[0m[38;2;148;128;130m█[0m[38;2;147;127;129m█[0m[38;2;144;126;125m█[0m[38;2;93;81;81m█[0m[38;2;135;129;129m█[0m[38;2;199;199;201m█[0m[38;2;196;196;202m█[0m[38;2;191;190;196m█[0m[38;2;190;189;195m█[0m[38;2;192;191;197m█[0m[38;2;186;185;188m█[0m[38;2;79;74;73m█[0m[38;2;142;139;139m█[0m");
		$display("[38;2;196;195;201m█[0m[38;2;199;197;202m█[0m[38;2;105;99;101m█[0m[38;2;107;104;104m█[0m[38;2;194;196;198m█[0m[38;2;192;190;197m█[0m[38;2;193;192;198m█[0m[38;2;194;193;199m█[0m[38;2;196;195;201m█[0m[38;2;198;197;203m█[0m[38;2;188;187;192m█[0m[38;2;86;80;81m█[0m[38;2;168;166;169m█[0m[38;2;198;197;202m█[0m[38;2;195;194;200m██[0m[38;2;194;193;199m█[0m[38;2;192;191;197m██[0m[38;2;200;199;205m█[0m[38;2;118;114;117m█[0m[38;2;144;140;142m█[0m[38;2;202;202;207m█[0m[38;2;191;188;191m█[0m[38;2;119;93;91m█[0m[38;2;184;176;180m█[0m[38;2;195;196;201m█[0m[38;2;200;199;204m█[0m[38;2;140;136;139m█[0m[38;2;95;86;89m█[0m[38;2;198;197;202m█[0m[38;2;192;191;197m█[0m[38;2;191;190;196m█[0m[38;2;194;193;199m█[0m[38;2;197;196;202m██[0m[38;2;202;201;205m█[0m[38;2;108;105;105m█[0m[38;2;116;107;106m█[0m[38;2;120;101;104m█[0m[38;2;110;90;90m█[0m[38;2;164;151;149m█[0m[38;2;202;193;191m█[0m[38;2;103;95;93m█[0m[38;2;157;148;147m█[0m[38;2;223;216;214m█[0m[38;2;212;203;203m█[0m[38;2;211;201;201m█[0m[38;2;210;198;198m█[0m[38;2;209;199;198m█[0m[38;2;178;169;167m█[0m[38;2;85;76;74m█[0m[38;2;192;181;181m█[0m[38;2;207;196;197m█[0m[38;2;212;202;202m█[0m[38;2;218;210;208m█[0m[38;2;222;214;211m█[0m[38;2;88;81;79m█[0m[38;2;175;167;165m█[0m[38;2;218;212;209m█[0m[38;2;190;178;177m█[0m[38;2;144;128;127m█[0m[38;2;106;89;88m█[0m[38;2;119;104;103m█[0m[38;2;100;95;95m█[0m[38;2;160;158;159m█[0m[38;2;146;134;136m█[0m[38;2;196;195;199m█[0m[38;2;184;180;186m█[0m[38;2;163;157;160m█[0m[38;2;198;197;201m█[0m[38;2;201;199;205m█[0m[38;2;101;94;97m█[0m[38;2;140;137;139m█[0m[38;2;199;199;204m█[0m[38;2;193;192;198m██[0m[38;2;194;193;199m█[0m[38;2;196;195;201m█[0m[38;2;199;198;204m█[0m[38;2;170;169;172m█[0m[38;2;87;84;84m█[0m[38;2;192;191;194m█[0m[38;2;197;197;202m█[0m[38;2;200;200;206m█[0m[38;2;202;202;208m█[0m[38;2;197;195;201m█[0m[38;2;190;185;191m█[0m[38;2;190;185;192m█[0m[38;2;201;198;203m█[0m[38;2;110;107;108m█[0m[38;2;137;135;136m█[0m[38;2;200;199;203m█[0m[38;2;194;193;199m██[0m[38;2;192;191;197m█[0m[38;2;195;194;200m█[0m[38;2;177;176;178m█[0m[38;2;71;66;65m█[0m[38;2;154;153;154m█[0m");
        $display("********************************************************");     
        $display("                     FAIL!                              ");
        $display("*                 Wrong answer                         *");
        $display("********************************************************");
        repeat(2) @(negedge clk);
        $finish;
    end
    @(negedge clk);
end endtask

task YOU_PASS_task; begin
	$display("[38;2;245;199;150m█[0m[38;2;247;201;152m█[0m[38;2;246;200;152m█[0m[38;2;244;199;153m█[0m[38;2;232;189;144m█[0m[38;2;226;183;138m█[0m[38;2;227;183;136m█[0m[38;2;235;191;142m█[0m[38;2;243;200;151m█[0m[38;2;247;205;157m██[0m[38;2;246;204;156m█[0m[38;2;245;203;155m█[0m[38;2;244;200;153m█[0m[38;2;245;201;154m█[0m[38;2;245;203;155m█[0m[38;2;246;204;156m█[0m[38;2;246;204;155m█[0m[38;2;245;203;156m█[0m[38;2;245;202;159m█[0m[38;2;246;204;162m█[0m[38;2;248;206;164m██[0m[38;2;247;205;163m█[0m[38;2;245;204;160m██[0m[38;2;247;206;162m██[0m[38;2;243;202;157m█[0m[38;2;230;189;144m█[0m[38;2;238;197;151m█[0m[38;2;242;200;157m█[0m[38;2;245;204;163m█[0m[38;2;246;208;167m█[0m[38;2;247;210;168m█[0m[38;2;246;208;164m█[0m[38;2;247;205;161m█[0m[38;2;248;205;161m█[0m[38;2;247;206;164m█[0m[38;2;247;209;169m█[0m[38;2;247;209;170m█[0m[38;2;246;208;169m█[0m[38;2;245;208;166m█[0m[38;2;245;207;163m█[0m[38;2;248;208;165m█[0m[38;2;221;195;163m█[0m[38;2;167;158;147m█[0m[38;2;221;187;153m█[0m[38;2;86;53;49m█[0m[38;2;205;159;164m█[0m[38;2;249;199;207m█[0m[38;2;246;195;205m█[0m[38;2;244;199;203m█[0m[38;2;248;232;207m█[0m[38;2;254;245;210m█[0m[38;2;246;236;205m█[0m[38;2;109;90;81m█[0m[38;2;113;83;67m█[0m[38;2;238;200;159m█[0m[38;2;254;215;169m█[0m[38;2;192;156;129m█[0m[38;2;95;61;61m█[0m[38;2;222;178;185m█[0m[38;2;248;199;208m█[0m[38;2;245;195;205m█[0m[38;2;244;197;204m█[0m[38;2;246;221;205m█[0m[38;2;251;240;208m█[0m[38;2;253;243;210m█[0m[38;2;255;248;216m█[0m[38;2;198;188;163m█[0m[38;2;100;81;66m█[0m[38;2;155;126;102m█[0m[38;2;242;204;160m█[0m[38;2;247;205;161m█[0m[38;2;246;204;160m█[0m[38;2;243;201;159m█[0m[38;2;233;191;149m█[0m[38;2;228;186;143m█[0m[38;2;239;197;151m█[0m[38;2;247;205;157m█[0m[38;2;246;204;156m█[0m[38;2;240;198;151m█[0m[38;2;228;186;141m█[0m[38;2;223;180;137m█[0m[38;2;235;192;147m█[0m[38;2;245;203;155m█[0m[38;2;243;201;153m█[0m[38;2;241;199;151m█[0m[38;2;239;197;149m██[0m[38;2;234;192;144m█[0m[38;2;228;186;138m█[0m[38;2;226;183;134m█[0m[38;2;237;193;144m█[0m[38;2;245;201;151m█[0m[38;2;246;200;150m█[0m[38;2;244;198;148m█[0m[38;2;244;197;145m██[0m");
	$display("[38;2;246;200;151m█[0m[38;2;247;201;151m█[0m[38;2;246;200;151m█[0m[38;2;245;200;151m█[0m[38;2;246;202;154m█[0m[38;2;246;202;155m█[0m[38;2;241;198;150m█[0m[38;2;232;188;141m█[0m[38;2;227;182;136m█[0m[38;2;228;184;141m█[0m[38;2;236;192;148m█[0m[38;2;243;201;153m█[0m[38;2;245;203;155m█[0m[38;2;247;204;156m█[0m[38;2;246;203;155m█[0m[38;2;245;202;154m█[0m[38;2;246;204;156m█[0m[38;2;246;204;157m█[0m[38;2;245;203;157m█[0m[38;2;247;204;160m█[0m[38;2;247;205;162m█[0m[38;2;246;205;161m█[0m[38;2;245;204;159m█[0m[38;2;246;204;159m█[0m[38;2;246;205;159m█[0m[38;2;248;206;162m█[0m[38;2;248;206;164m██[0m[38;2;247;206;163m██[0m[38;2;240;199;156m█[0m[38;2;241;199;157m█[0m[38;2;245;204;163m█[0m[38;2;246;207;167m█[0m[38;2;246;208;166m█[0m[38;2;247;208;165m█[0m[38;2;248;206;163m██[0m[38;2;247;208;164m█[0m[38;2;248;210;168m█[0m[38;2;248;210;169m█[0m[38;2;247;209;167m█[0m[38;2;246;207;166m█[0m[38;2;246;208;165m█[0m[38;2;249;210;167m█[0m[38;2;187;173;157m█[0m[38;2;185;171;155m█[0m[38;2;194;159;129m█[0m[38;2;95;66;64m█[0m[38;2;238;191;197m█[0m[38;2;246;196;206m█[0m[38;2;245;196;204m█[0m[38;2;248;223;207m█[0m[38;2;252;244;208m█[0m[38;2;251;243;209m█[0m[38;2;128;112;95m█[0m[38;2;98;66;57m█[0m[38;2;233;198;161m█[0m[38;2;252;214;169m█[0m[38;2;224;190;156m█[0m[38;2;94;63;59m█[0m[38;2;196;153;159m█[0m[38;2;252;201;210m█[0m[38;2;245;194;204m█[0m[38;2;245;205;203m█[0m[38;2;249;230;205m█[0m[38;2;251;241;208m█[0m[38;2;255;247;213m█[0m[38;2;241;231;201m█[0m[38;2;140;126;106m█[0m[38;2;102;80;60m█[0m[38;2;200;165;130m█[0m[38;2;252;210;167m█[0m[38;2;249;207;163m█[0m[38;2;244;202;160m█[0m[38;2;236;194;152m█[0m[38;2;234;192;150m█[0m[38;2;241;199;157m█[0m[38;2;246;205;162m█[0m[38;2;246;204;160m█[0m[38;2;238;197;153m█[0m[38;2;228;187;143m█[0m[38;2;230;188;143m█[0m[38;2;239;197;154m█[0m[38;2;244;203;158m█[0m[38;2;242;201;153m█[0m[38;2;242;199;152m█[0m[38;2;242;201;152m█[0m[38;2;238;197;149m█[0m[38;2;235;193;145m█[0m[38;2;235;192;144m█[0m[38;2;237;195;147m█[0m[38;2;243;202;153m█[0m[38;2;247;203;156m█[0m[38;2;247;202;155m█[0m[38;2;246;202;154m█[0m[38;2;245;199;150m█[0m[38;2;246;198;148m█[0m[38;2;246;198;149m█[0m[38;2;245;197;148m█[0m");
	$display("[38;2;247;201;151m██[0m[38;2;246;200;150m█[0m[38;2;245;199;150m█[0m[38;2;245;200;151m█[0m[38;2;245;201;152m█[0m[38;2;245;202;154m█[0m[38;2;246;202;155m█[0m[38;2;246;201;155m█[0m[38;2;241;198;152m█[0m[38;2;235;192;146m█[0m[38;2;230;188;140m██[0m[38;2;236;193;147m█[0m[38;2;242;200;154m█[0m[38;2;246;203;157m█[0m[38;2;246;204;158m█[0m[38;2;246;204;159m█[0m[38;2;246;205;159m█[0m[38;2;247;206;161m█[0m[38;2;248;207;162m█[0m[38;2;247;206;161m█[0m[38;2;247;206;160m██[0m[38;2;247;206;162m█[0m[38;2;247;208;164m█[0m[38;2;248;206;164m█[0m[38;2;249;206;165m█[0m[38;2;247;207;164m█[0m[38;2;247;208;165m█[0m[38;2;248;208;166m█[0m[38;2;247;206;165m█[0m[38;2;247;207;165m█[0m[38;2;249;209;168m█[0m[38;2;249;209;169m█[0m[38;2;249;208;167m█[0m[38;2;249;210;166m█[0m[38;2;247;209;167m█[0m[38;2;244;208;168m█[0m[38;2;243;209;171m█[0m[38;2;245;210;170m█[0m[38;2;252;214;172m█[0m[38;2;250;212;172m█[0m[38;2;247;209;169m█[0m[38;2;218;190;159m█[0m[38;2;174;160;147m█[0m[38;2;205;180;155m█[0m[38;2;152;120;97m█[0m[38;2;131;98;99m█[0m[38;2;250;201;208m█[0m[38;2;245;201;204m█[0m[38;2;248;225;206m█[0m[38;2;251;242;208m█[0m[38;2;252;245;210m█[0m[38;2;175;161;139m█[0m[38;2;69;42;35m█[0m[38;2;219;184;152m█[0m[38;2;255;219;180m█[0m[38;2;252;217;177m█[0m[38;2;122;93;80m█[0m[38;2;150;111;118m█[0m[38;2;252;202;212m█[0m[38;2;244;197;204m█[0m[38;2;246;216;203m█[0m[38;2;250;239;207m█[0m[38;2;251;242;207m█[0m[38;2;255;248;214m█[0m[38;2;212;201;176m█[0m[38;2;98;77;62m█[0m[38;2;135;105;82m█[0m[38;2;238;201;162m█[0m[38;2;253;214;170m█[0m[38;2;246;205;163m█[0m[38;2;240;199;157m█[0m[38;2;238;196;155m█[0m[38;2;243;201;161m█[0m[38;2;248;206;164m█[0m[38;2;246;204;162m█[0m[38;2;235;193;151m█[0m[38;2;231;190;148m█[0m[38;2;236;194;153m█[0m[38;2;243;201;160m█[0m[38;2;246;205;162m█[0m[38;2;245;204;160m█[0m[38;2;243;202;157m█[0m[38;2;242;201;156m█[0m[38;2;239;198;151m█[0m[38;2;239;198;150m█[0m[38;2;242;200;152m█[0m[38;2;245;204;157m█[0m[38;2;247;206;159m█[0m[38;2;247;205;159m█[0m[38;2;247;204;158m█[0m[38;2;245;202;155m█[0m[38;2;245;201;154m█[0m[38;2;245;201;153m█[0m[38;2;242;197;148m█[0m[38;2;241;194;145m█[0m[38;2;241;194;144m█[0m[38;2;241;194;146m█[0m");
	$display("[38;2;246;200;150m█[0m[38;2;245;200;151m█[0m[38;2;245;199;150m█[0m[38;2;245;200;150m█[0m[38;2;245;200;152m█[0m[38;2;245;201;152m█[0m[38;2;246;202;153m█[0m[38;2;246;202;154m█[0m[38;2;246;203;155m█[0m[38;2;246;204;157m█[0m[38;2;247;205;158m██[0m[38;2;245;203;156m█[0m[38;2;240;198;153m█[0m[38;2;235;193;149m█[0m[38;2;235;194;149m█[0m[38;2;238;196;151m█[0m[38;2;242;201;155m█[0m[38;2;247;206;160m█[0m[38;2;248;207;163m█[0m[38;2;248;207;164m███[0m[38;2;247;207;164m█[0m[38;2;247;206;164m█[0m[38;2;247;208;165m█[0m[38;2;248;207;164m█[0m[38;2;248;207;165m█[0m[38;2;247;208;165m█[0m[38;2;248;209;166m█[0m[38;2;250;211;167m█[0m[38;2;250;211;169m█[0m[38;2;245;208;168m█[0m[38;2;238;204;168m█[0m[38;2;228;197;169m█[0m[38;2;212;187;161m█[0m[38;2;197;173;149m█[0m[38;2;183;157;134m█[0m[38;2;170;144;121m█[0m[38;2;163;137;119m█[0m[38;2;158;132;110m█[0m[38;2;158;131;106m█[0m[38;2;151;125;104m█[0m[38;2;148;122;103m█[0m[38;2;147;123;103m█[0m[38;2;151;126;109m█[0m[38;2;153;131;109m█[0m[38;2;136;116;99m█[0m[38;2;202;180;162m█[0m[38;2;252;231;211m█[0m[38;2;250;236;208m█[0m[38;2;251;242;208m█[0m[38;2;254;245;211m█[0m[38;2;190;180;152m█[0m[38;2;113;96;80m█[0m[38;2;114;90;77m█[0m[38;2;148;122;100m█[0m[38;2;152;124;102m█[0m[38;2;144;118;99m█[0m[38;2;104;74;73m█[0m[38;2;238;192;197m█[0m[38;2;247;208;205m█[0m[38;2;249;229;205m█[0m[38;2;252;241;209m█[0m[38;2;251;241;207m█[0m[38;2;255;247;213m█[0m[38;2;191;179;154m█[0m[38;2;85;61;50m█[0m[38;2;178;144;117m█[0m[38;2;252;214;172m█[0m[38;2;246;208;166m█[0m[38;2;242;204;161m█[0m[38;2;242;204;162m█[0m[38;2;246;207;166m█[0m[38;2;248;206;165m█[0m[38;2;244;202;161m█[0m[38;2;237;195;153m██[0m[38;2;240;198;156m█[0m[38;2;246;204;162m██[0m[38;2;244;202;160m██[0m[38;2;243;202;159m█[0m[38;2;244;203;160m█[0m[38;2;245;204;159m█[0m[38;2;245;204;155m█[0m[38;2;246;204;156m██[0m[38;2;246;202;156m█[0m[38;2;244;201;155m█[0m[38;2;241;198;152m█[0m[38;2;239;195;150m█[0m[38;2;237;192;146m█[0m[38;2;237;192;145m█[0m[38;2;240;195;148m█[0m[38;2;242;199;150m█[0m[38;2;247;203;153m█[0m[38;2;248;202;152m█[0m[38;2;248;201;153m█[0m");
	$display("[38;2;246;200;151m█[0m[38;2;246;202;153m█[0m[38;2;245;202;153m██[0m[38;2;245;202;154m█[0m[38;2;246;203;156m█[0m[38;2;246;203;157m██[0m[38;2;246;204;158m█[0m[38;2;247;204;160m█[0m[38;2;247;205;160m███[0m[38;2;247;207;162m█[0m[38;2;247;206;162m█[0m[38;2;246;205;162m█[0m[38;2;244;203;159m█[0m[38;2;240;199;154m█[0m[38;2;239;197;153m█[0m[38;2;241;200;157m█[0m[38;2;244;203;159m█[0m[38;2;247;205;162m█[0m[38;2;249;207;165m█[0m[38;2;248;208;165m█[0m[38;2;248;206;164m█[0m[38;2;247;207;165m█[0m[38;2;248;209;166m█[0m[38;2;251;211;167m█[0m[38;2;248;209;168m█[0m[38;2;237;203;167m█[0m[38;2;223;195;164m█[0m[38;2;210;187;164m█[0m[38;2;193;172;151m█[0m[38;2;166;144;125m█[0m[38;2;140;119;101m█[0m[38;2;135;113;96m█[0m[38;2;148;126;108m█[0m[38;2;167;149;128m█[0m[38;2;184;168;144m█[0m[38;2;201;186;161m█[0m[38;2;215;203;176m█[0m[38;2;225;215;186m█[0m[38;2;235;225;195m█[0m[38;2;242;232;201m█[0m[38;2;247;237;205m█[0m[38;2;250;240;208m█[0m[38;2;252;242;209m█[0m[38;2;255;246;212m█[0m[38;2;254;244;211m█[0m[38;2;251;241;208m██[0m[38;2;251;240;208m█[0m[38;2;251;241;208m█[0m[38;2;249;239;206m██[0m[38;2;250;240;206m█[0m[38;2;242;232;201m█[0m[38;2;232;221;192m█[0m[38;2;217;205;177m█[0m[38;2;234;220;193m█[0m[38;2;252;236;209m█[0m[38;2;251;240;207m█[0m[38;2;251;242;207m█[0m[38;2;251;240;208m█[0m[38;2;254;245;212m█[0m[38;2;208;198;170m█[0m[38;2;92;69;55m█[0m[38;2;205;169;137m█[0m[38;2;255;217;173m█[0m[38;2;251;211;168m█[0m[38;2;251;211;169m█[0m[38;2;251;212;170m█[0m[38;2;249;210;169m█[0m[38;2;244;206;164m█[0m[38;2;241;200;158m██[0m[38;2;244;202;160m█[0m[38;2;247;205;163m██[0m[38;2;246;204;162m█[0m[38;2;246;205;162m█[0m[38;2;247;205;162m█[0m[38;2;246;205;162m█[0m[38;2;247;205;163m██[0m[38;2;246;205;160m█[0m[38;2;245;203;154m█[0m[38;2;243;202;153m█[0m[38;2;239;197;149m█[0m[38;2;236;192;145m██[0m[38;2;239;196;148m█[0m[38;2;244;200;153m█[0m[38;2;248;204;157m█[0m[38;2;249;205;158m█[0m[38;2;244;201;155m█[0m[38;2;234;190;148m█[0m[38;2;219;176;136m█[0m[38;2;201;160;122m█[0m[38;2;187;147;111m█[0m");
	$display("[38;2;245;200;151m█[0m[38;2;246;202;153m███[0m[38;2;245;203;154m█[0m[38;2;246;204;156m█[0m[38;2;246;204;157m█[0m[38;2;247;204;158m█[0m[38;2;246;204;159m█[0m[38;2;246;205;160m█[0m[38;2;247;206;161m█[0m[38;2;247;206;162m█[0m[38;2;248;207;163m█[0m[38;2;246;204;160m██[0m[38;2;247;205;163m█[0m[38;2;248;206;164m█[0m[38;2;248;207;164m█[0m[38;2;248;206;164m█[0m[38;2;246;204;162m█[0m[38;2;244;202;160m██[0m[38;2;246;204;162m█[0m[38;2;248;206;164m█[0m[38;2;249;209;167m█[0m[38;2;249;209;168m█[0m[38;2;234;200;161m█[0m[38;2;214;189;163m█[0m[38;2;207;183;158m█[0m[38;2;197;173;147m█[0m[38;2;171;145;126m█[0m[38;2;152;125;106m█[0m[38;2;152;131;111m█[0m[38;2;180;164;143m█[0m[38;2;215;204;175m█[0m[38;2;241;231;199m█[0m[38;2;253;243;210m█[0m[38;2;255;247;214m██[0m[38;2;255;246;213m██[0m[38;2;255;245;212m███[0m[38;2;254;243;211m█[0m[38;2;252;241;209m█[0m[38;2;251;240;208m████████[0m[38;2;252;241;209m███[0m[38;2;253;242;210m█[0m[38;2;255;244;211m█[0m[38;2;254;243;210m█[0m[38;2;251;241;208m█[0m[38;2;251;240;208m███[0m[38;2;252;242;210m█[0m[38;2;228;217;187m█[0m[38;2;223;206;175m█[0m[38;2;255;235;199m█[0m[38;2;216;189;157m█[0m[38;2;181;151;123m█[0m[38;2;185;153;122m█[0m[38;2;203;168;133m█[0m[38;2;229;192;153m█[0m[38;2;245;208;166m█[0m[38;2;250;212;169m█[0m[38;2;249;210;167m█[0m[38;2;248;206;164m█[0m[38;2;247;205;164m██[0m[38;2;247;205;162m█[0m[38;2;246;206;162m█[0m[38;2;247;207;164m██[0m[38;2;248;206;164m█[0m[38;2;246;204;162m█[0m[38;2;246;205;160m█[0m[38;2;246;205;157m█[0m[38;2;245;205;156m█[0m[38;2;246;204;156m█[0m[38;2;247;203;156m█[0m[38;2;242;199;154m█[0m[38;2;232;189;145m█[0m[38;2;216;176;133m█[0m[38;2;203;162;123m█[0m[38;2;193;150;115m█[0m[38;2;185;144;110m█[0m[38;2;189;150;112m█[0m[38;2;203;164;124m█[0m[38;2;219;178;137m█[0m[38;2;232;190;147m█[0m");
	$display("[38;2;245;203;155m██[0m[38;2;246;204;156m█[0m[38;2;245;203;155m███[0m[38;2;246;204;156m██[0m[38;2;246;203;156m█[0m[38;2;246;204;156m█[0m[38;2;246;204;157m█[0m[38;2;247;206;162m██[0m[38;2;247;204;161m█[0m[38;2;246;204;160m█[0m[38;2;247;206;162m██[0m[38;2;248;206;163m█[0m[38;2;248;206;164m█[0m[38;2;247;205;164m█[0m[38;2;247;206;164m█[0m[38;2;248;206;164m█[0m[38;2;250;210;166m█[0m[38;2;244;209;169m█[0m[38;2;218;194;167m█[0m[38;2;198;181;159m█[0m[38;2;203;182;157m█[0m[38;2;191;165;142m█[0m[38;2;150;122;104m█[0m[38;2;131;106;89m█[0m[38;2;166;148;126m█[0m[38;2;218;206;179m█[0m[38;2;249;240;208m█[0m[38;2;255;247;215m█[0m[38;2;255;244;212m█[0m[38;2;252;242;209m█[0m[38;2;253;243;210m█[0m[38;2;255;246;213m█[0m[38;2;255;245;213m█[0m[38;2;250;238;207m█[0m[38;2;239;228;197m█[0m[38;2;230;218;187m█[0m[38;2;223;211;180m█[0m[38;2;222;211;179m█[0m[38;2;230;219;187m█[0m[38;2;246;236;204m█[0m[38;2;251;240;208m███████████████[0m[38;2;252;241;208m██[0m[38;2;251;240;208m██[0m[38;2;253;243;210m█[0m[38;2;254;244;211m█[0m[38;2;251;241;209m█[0m[38;2;247;237;206m█[0m[38;2;234;224;195m█[0m[38;2;211;200;173m█[0m[38;2;179;164;141m█[0m[38;2;151;130;110m█[0m[38;2;145;118;97m█[0m[38;2;175;143;113m█[0m[38;2;221;185;147m█[0m[38;2;249;211;169m█[0m[38;2;252;212;170m█[0m[38;2;249;207;165m█[0m[38;2;248;206;164m█[0m[38;2;247;207;164m█[0m[38;2;247;209;166m█[0m[38;2;248;208;165m█[0m[38;2;249;208;165m█[0m[38;2;248;206;164m█[0m[38;2;243;203;161m█[0m[38;2;233;195;154m█[0m[38;2;221;182;141m█[0m[38;2;207;169;128m█[0m[38;2;196;156;120m█[0m[38;2;196;155;119m█[0m[38;2;201;162;125m█[0m[38;2;213;175;134m█[0m[38;2;225;185;141m█[0m[38;2;234;191;149m█[0m[38;2;233;192;151m█[0m[38;2;223;182;139m█[0m[38;2;207;165;128m█[0m[38;2;188;149;117m█[0m[38;2;171;134;106m█[0m");
	$display("[38;2;243;201;153m█[0m[38;2;242;201;153m█[0m[38;2;245;202;155m█[0m[38;2;245;202;157m█[0m[38;2;246;204;157m█[0m[38;2;245;203;155m█[0m[38;2;245;202;154m█[0m[38;2;245;201;154m█[0m[38;2;246;202;155m█[0m[38;2;245;202;156m█[0m[38;2;246;204;160m█[0m[38;2;247;206;162m█████[0m[38;2;248;207;163m█[0m[38;2;248;206;163m█[0m[38;2;249;206;164m█[0m[38;2;248;207;166m█[0m[38;2;249;209;167m█[0m[38;2;245;207;166m█[0m[38;2;218;190;158m█[0m[38;2;198;179;155m█[0m[38;2;210;188;165m█[0m[38;2;193;165;138m█[0m[38;2;137;112;93m█[0m[38;2;134;114;97m█[0m[38;2;191;178;156m█[0m[38;2;243;233;202m█[0m[38;2;255;248;215m█[0m[38;2;255;245;211m█[0m[38;2;251;241;208m█[0m[38;2;251;240;208m█[0m[38;2;255;244;211m█[0m[38;2;255;245;212m█[0m[38;2;232;222;190m█[0m[38;2;192;180;155m█[0m[38;2;162;149;127m█[0m[38;2;159;145;123m█[0m[38;2;169;155;133m█[0m[38;2;182;168;144m█[0m[38;2;190;176;151m█[0m[38;2;193;180;154m█[0m[38;2;196;184;158m█[0m[38;2;225;213;185m█[0m[38;2;253;242;210m█[0m[38;2;251;240;208m█████████████[0m[38;2;250;239;207m█[0m[38;2;245;235;202m█[0m[38;2;244;234;201m█[0m[38;2;248;238;204m█[0m[38;2;253;243;209m█[0m[38;2;255;246;213m█[0m[38;2;255;245;213m█[0m[38;2;253;242;210m█[0m[38;2;252;241;209m█[0m[38;2;253;242;209m█[0m[38;2;255;245;212m█[0m[38;2;255;247;214m█[0m[38;2;254;244;212m█[0m[38;2;233;221;193m█[0m[38;2;188;174;153m█[0m[38;2;144;124;107m█[0m[38;2;137;111;91m█[0m[38;2;187;153;122m█[0m[38;2;239;201;161m█[0m[38;2;253;215;171m█[0m[38;2;247;207;162m█[0m[38;2;240;199;156m█[0m[38;2;233;191;151m█[0m[38;2;225;183;143m█[0m[38;2;219;177;139m█[0m[38;2;215;175;139m█[0m[38;2;214;177;141m█[0m[38;2;221;183;144m█[0m[38;2;228;186;144m█[0m[38;2;230;187;145m█[0m[38;2;225;184;142m█[0m[38;2;213;173;134m█[0m[38;2;198;159;123m█[0m[38;2;188;149;116m█[0m[38;2;178;140;110m█[0m[38;2;171;135;106m█[0m[38;2;174;137;106m█[0m[38;2;183;144;112m█[0m[38;2;195;156;123m█[0m[38;2;207;168;133m█[0m");
	$display("[38;2;243;201;153m█[0m[38;2;242;200;152m█[0m[38;2;244;201;154m█[0m[38;2;244;202;154m█[0m[38;2;245;203;156m█[0m[38;2;245;203;157m█[0m[38;2;245;202;156m█[0m[38;2;246;202;157m█[0m[38;2;246;203;158m█[0m[38;2;246;204;160m█[0m[38;2;246;205;161m█[0m[38;2;247;205;161m██[0m[38;2;247;205;160m█[0m[38;2;246;204;159m█[0m[38;2;247;205;162m█[0m[38;2;248;206;164m█[0m[38;2;249;206;165m█[0m[38;2;250;207;165m█[0m[38;2;250;208;165m█[0m[38;2;225;195;162m█[0m[38;2;199;178;152m█[0m[38;2;221;194;163m█[0m[38;2;212;177;145m█[0m[38;2;138;107;86m█[0m[38;2;135;114;97m█[0m[38;2;207;195;170m█[0m[38;2;253;243;212m█[0m[38;2;255;247;213m█[0m[38;2;252;242;209m█[0m[38;2;251;240;208m██[0m[38;2;253;243;209m█[0m[38;2;255;245;212m█[0m[38;2;216;205;178m█[0m[38;2;164;150;130m█[0m[38;2;167;153;130m█[0m[38;2;200;188;162m█[0m[38;2;229;218;188m█[0m[38;2;247;236;205m█[0m[38;2;254;243;212m█[0m[38;2;255;246;213m███[0m[38;2;255;245;212m█[0m[38;2;253;242;209m█[0m[38;2;251;240;208m█████████████[0m[38;2;252;242;210m█[0m[38;2;224;213;182m█[0m[38;2;196;184;160m█[0m[38;2;187;175;152m█[0m[38;2;176;163;140m█[0m[38;2;170;157;134m█[0m[38;2;175;162;138m█[0m[38;2;201;188;161m█[0m[38;2;236;226;195m█[0m[38;2;255;247;214m█[0m[38;2;254;244;211m█[0m[38;2;251;240;208m███[0m[38;2;253;242;210m█[0m[38;2;255;247;213m█[0m[38;2;255;245;213m█[0m[38;2;223;213;185m█[0m[38;2;163;146;129m█[0m[38;2;129;105;89m█[0m[38;2;159;129;103m█[0m[38;2;220;181;146m█[0m[38;2;242;201;162m█[0m[38;2;238;196;155m█[0m[38;2;237;195;153m█[0m[38;2;236;194;153m█[0m[38;2;234;191;153m█[0m[38;2;229;186;148m█[0m[38;2;221;179;140m█[0m[38;2;219;177;139m█[0m[38;2;217;175;137m█[0m[38;2;215;174;136m█[0m[38;2;220;180;143m█[0m[38;2;226;185;148m█[0m[38;2;234;194;155m█[0m[38;2;241;201;159m█[0m[38;2;245;205;161m█[0m[38;2;248;206;158m█[0m[38;2;249;207;155m█[0m[38;2;250;207;158m█[0m[38;2;251;206;159m█[0m");
	$display("[38;2;246;203;155m█[0m[38;2;247;204;156m█[0m[38;2;246;203;155m██[0m[38;2;246;203;157m█[0m[38;2;246;205;159m██[0m[38;2;246;204;157m█[0m[38;2;246;204;159m█[0m[38;2;246;205;161m███[0m[38;2;247;205;162m█[0m[38;2;247;205;161m█[0m[38;2;247;206;162m█[0m[38;2;247;206;164m█[0m[38;2;248;206;165m█[0m[38;2;250;208;165m█[0m[38;2;243;205;167m█[0m[38;2;202;179;155m█[0m[38;2;209;187;161m█[0m[38;2;235;199;162m█[0m[38;2;155;123;97m█[0m[38;2;108;86;72m█[0m[38;2;194;183;157m█[0m[38;2;255;246;213m██[0m[38;2;251;240;208m███[0m[38;2;251;240;207m█[0m[38;2;255;246;212m█[0m[38;2;233;221;194m█[0m[38;2;164;150;128m█[0m[38;2;172;158;136m█[0m[38;2;228;216;188m█[0m[38;2;255;245;213m█[0m[38;2;255;246;213m█[0m[38;2;253;242;210m█[0m[38;2;252;241;208m█[0m[38;2;251;240;208m████████████████████[0m[38;2;252;241;209m█[0m[38;2;253;243;210m██[0m[38;2;251;240;208m█[0m[38;2;243;232;200m█[0m[38;2;224;212;183m█[0m[38;2;191;179;153m█[0m[38;2;159;145;125m█[0m[38;2;164;150;125m█[0m[38;2;222;210;179m█[0m[38;2;255;247;214m█[0m[38;2;252;242;208m█[0m[38;2;251;240;208m████[0m[38;2;254;244;210m█[0m[38;2;255;248;215m█[0m[38;2;241;232;201m█[0m[38;2;180;167;145m█[0m[38;2;128;105;87m█[0m[38;2;167;135;110m█[0m[38;2;229;191;150m█[0m[38;2;242;199;157m█[0m[38;2;237;195;153m█[0m[38;2;240;198;158m█[0m[38;2;243;201;161m█[0m[38;2;246;205;161m█[0m[38;2;248;207;163m█[0m[38;2;249;208;164m██[0m[38;2;248;207;163m█[0m[38;2;248;207;161m█[0m[38;2;247;205;161m█[0m[38;2;246;205;161m█[0m[38;2;245;204;160m█[0m[38;2;245;204;159m█[0m[38;2;245;203;156m█[0m[38;2;246;203;155m██[0m");
	$display("[38;2;239;195;148m█[0m[38;2;241;198;151m█[0m[38;2;243;200;153m█[0m[38;2;244;201;153m█[0m[38;2;245;201;156m█[0m[38;2;245;202;157m█[0m[38;2;246;204;157m█[0m[38;2;247;205;157m█[0m[38;2;247;205;158m█[0m[38;2;247;206;161m█[0m[38;2;248;207;163m█[0m[38;2;248;207;164m█[0m[38;2;248;206;164m█[0m[38;2;248;206;163m█[0m[38;2;248;206;164m█[0m[38;2;247;207;165m█[0m[38;2;250;210;168m█[0m[38;2;235;201;167m█[0m[38;2;184;168;153m█[0m[38;2;225;199;169m█[0m[38;2;215;178;146m█[0m[38;2;104;74;58m█[0m[38;2;133;117;102m█[0m[38;2;238;228;200m█[0m[38;2;255;247;215m█[0m[38;2;251;240;208m█████[0m[38;2;255;246;212m█[0m[38;2;211;200;172m█[0m[38;2;154;140;120m█[0m[38;2;222;209;182m█[0m[38;2;255;247;214m█[0m[38;2;254;243;210m█[0m[38;2;251;240;208m████████████████████████████[0m[38;2;252;241;209m█[0m[38;2;254;243;211m█[0m[38;2;255;246;214m█[0m[38;2;254;243;212m█[0m[38;2;222;210;182m█[0m[38;2;160;147;124m█[0m[38;2;171;158;134m█[0m[38;2;247;237;205m█[0m[38;2;254;243;211m█[0m[38;2;251;240;208m█████[0m[38;2;253;242;209m█[0m[38;2;255;248;214m█[0m[38;2;243;235;202m█[0m[38;2;172;155;138m█[0m[38;2;120;93;74m█[0m[38;2;190;154;117m█[0m[38;2;251;211;166m█[0m[38;2;249;207;163m█[0m[38;2;245;204;160m█[0m[38;2;245;204;161m█[0m[38;2;245;204;160m█[0m[38;2;245;204;161m█[0m[38;2;246;205;161m█[0m[38;2;245;204;160m█[0m[38;2;243;202;158m█[0m[38;2;243;202;157m█[0m[38;2;244;203;157m█[0m[38;2;243;203;156m█[0m[38;2;243;203;155m█[0m[38;2;245;202;156m█[0m[38;2;245;204;155m█[0m[38;2;246;204;156m█[0m");
	$display("[38;2;233;190;145m█[0m[38;2;235;192;147m█[0m[38;2;234;194;149m█[0m[38;2;234;192;149m█[0m[38;2;234;191;147m█[0m[38;2;235;192;147m█[0m[38;2;236;193;149m█[0m[38;2;237;195;150m█[0m[38;2;239;197;152m█[0m[38;2;243;202;156m█[0m[38;2;244;202;158m█[0m[38;2;246;204;161m█[0m[38;2;246;204;162m█[0m[38;2;246;204;163m█[0m[38;2;247;205;164m█[0m[38;2;250;209;168m█[0m[38;2;234;200;169m█[0m[38;2;175;164;150m█[0m[38;2;230;202;172m█[0m[38;2;189;155;126m█[0m[38;2;85;60;48m█[0m[38;2;178;165;142m█[0m[38;2;255;247;215m█[0m[38;2;254;244;209m█[0m[38;2;251;240;208m█████[0m[38;2;254;244;212m█[0m[38;2;218;206;179m█[0m[38;2;163;150;127m█[0m[38;2;247;237;205m█[0m[38;2;255;245;212m█[0m[38;2;251;240;208m██████[0m[38;2;253;242;210m█[0m[38;2;255;244;211m█[0m[38;2;254;243;211m█[0m[38;2;252;241;209m█[0m[38;2;251;240;208m████████████████████████[0m[38;2;255;244;211m█[0m[38;2;255;246;214m█[0m[38;2;198;185;162m█[0m[38;2;145;132;109m█[0m[38;2;236;226;196m█[0m[38;2;254;244;212m█[0m[38;2;251;240;208m██████[0m[38;2;252;242;208m█[0m[38;2;255;249;216m█[0m[38;2;227;217;189m█[0m[38;2;132;111;95m█[0m[38;2;143;111;88m█[0m[38;2;238;200;160m█[0m[38;2;251;209;164m█[0m[38;2;245;207;163m█[0m[38;2;246;208;165m██[0m[38;2;247;208;165m█[0m[38;2;247;206;164m█[0m[38;2;245;204;160m█[0m[38;2;246;206;159m█[0m[38;2;247;206;160m█[0m[38;2;247;206;159m█[0m[38;2;245;203;155m████[0m");
	$display("[38;2;247;205;157m██[0m[38;2;247;205;158m█[0m[38;2;247;204;158m█[0m[38;2;246;204;158m█[0m[38;2;246;205;158m█[0m[38;2;245;205;158m█[0m[38;2;245;205;157m█[0m[38;2;245;204;157m█[0m[38;2;245;204;159m█[0m[38;2;246;204;161m█[0m[38;2;246;204;162m█[0m[38;2;246;205;162m█[0m[38;2;246;207;164m█[0m[38;2;248;209;169m█[0m[38;2;237;203;170m█[0m[38;2;171;158;146m█[0m[38;2;227;199;167m█[0m[38;2;181;146;121m█[0m[38;2;83;61;49m█[0m[38;2;204;193;167m█[0m[38;2;255;250;215m█[0m[38;2;252;241;208m█[0m[38;2;251;240;208m██████[0m[38;2;250;240;207m█[0m[38;2;178;165;140m█[0m[38;2;243;231;202m█[0m[38;2;253;244;209m█[0m[38;2;251;240;208m█████[0m[38;2;253;243;210m█[0m[38;2;255;246;214m█[0m[38;2;235;223;192m█[0m[38;2;218;206;176m█[0m[38;2;221;210;180m█[0m[38;2;247;236;205m█[0m[38;2;255;247;214m█[0m[38;2;251;241;208m█[0m[38;2;251;240;208m█████████████[0m[38;2;252;241;208m█[0m[38;2;253;242;210m█[0m[38;2;254;243;211m█[0m[38;2;253;243;210m█[0m[38;2;252;241;208m█[0m[38;2;251;240;208m█████[0m[38;2;251;240;207m█[0m[38;2;255;248;216m█[0m[38;2;210;199;172m█[0m[38;2;137;125;101m█[0m[38;2;244;235;203m█[0m[38;2;252;241;209m█[0m[38;2;251;240;208m███████[0m[38;2;255;244;212m█[0m[38;2;254;244;213m█[0m[38;2;169;152;134m█[0m[38;2;116;89;70m█[0m[38;2;226;190;150m█[0m[38;2;252;213;169m█[0m[38;2;246;207;165m█[0m[38;2;246;208;165m█[0m[38;2;247;208;165m█[0m[38;2;247;206;163m█[0m[38;2;245;205;159m█[0m[38;2;246;205;158m█[0m[38;2;246;205;159m█[0m[38;2;247;206;159m█[0m[38;2;247;205;157m█[0m[38;2;246;205;157m█[0m[38;2;245;204;155m█[0m[38;2;245;203;154m█[0m");
	$display("[38;2;240;198;150m█[0m[38;2;242;201;152m█[0m[38;2;244;202;153m█[0m[38;2;245;203;155m█[0m[38;2;246;204;157m█[0m[38;2;246;205;159m█[0m[38;2;246;205;160m██[0m[38;2;246;205;161m█[0m[38;2;246;204;162m███[0m[38;2;245;204;162m█[0m[38;2;245;206;163m█[0m[38;2;243;207;168m█[0m[38;2;175;161;146m█[0m[38;2;211;187;159m█[0m[38;2;186;155;124m█[0m[38;2;80;57;48m█[0m[38;2;211;199;173m█[0m[38;2;255;248;215m█[0m[38;2;251;240;208m███████[0m[38;2;252;241;208m█[0m[38;2;251;241;208m█[0m[38;2;248;238;205m█[0m[38;2;253;243;210m█[0m[38;2;251;241;208m███[0m[38;2;251;240;208m██[0m[38;2;252;243;210m█[0m[38;2;238;226;198m█[0m[38;2;142;126;109m█[0m[38;2;142;131;123m█[0m[38;2;173;165;160m█[0m[38;2;168;160;155m█[0m[38;2;118;103;92m█[0m[38;2;182;168;144m█[0m[38;2;251;242;210m█[0m[38;2;251;240;208m████████████[0m[38;2;255;246;212m█[0m[38;2;252;242;208m█[0m[38;2;231;220;188m█[0m[38;2;220;209;178m█[0m[38;2;229;217;186m█[0m[38;2;253;242;210m█[0m[38;2;255;246;213m█[0m[38;2;251;240;208m█████[0m[38;2;251;240;207m█[0m[38;2;255;249;216m█[0m[38;2;187;174;150m█[0m[38;2;170;156;130m█[0m[38;2;255;246;214m█[0m[38;2;251;240;208m████████[0m[38;2;252;241;208m█[0m[38;2;255;249;217m█[0m[38;2;190;175;154m█[0m[38;2;107;80;64m█[0m[38;2;225;190;152m█[0m[38;2;249;211;168m█[0m[38;2;247;205;163m██[0m[38;2;247;205;162m█[0m[38;2;246;206;160m█[0m[38;2;245;205;156m██[0m[38;2;246;206;158m█[0m[38;2;246;205;159m██[0m[38;2;246;206;158m█[0m[38;2;246;205;158m█[0m");
	$display("[38;2;244;202;156m█[0m[38;2;245;202;157m█[0m[38;2;245;203;157m█[0m[38;2;246;203;157m█[0m[38;2;246;203;158m██[0m[38;2;246;203;159m█[0m[38;2;246;203;160m█[0m[38;2;245;203;159m██[0m[38;2;245;203;161m█[0m[38;2;245;204;162m█[0m[38;2;245;205;163m█[0m[38;2;246;207;165m█[0m[38;2;192;173;150m█[0m[38;2;186;171;152m█[0m[38;2;215;180;147m█[0m[38;2;77;52;43m█[0m[38;2;192;177;158m█[0m[38;2;255;250;215m█[0m[38;2;251;240;208m██████[0m[38;2;251;242;207m██[0m[38;2;250;239;208m█[0m[38;2;250;233;210m█[0m[38;2;250;230;207m█[0m[38;2;249;229;206m█[0m[38;2;249;230;206m█[0m[38;2;248;230;206m█[0m[38;2;250;234;207m█[0m[38;2;251;241;208m█[0m[38;2;251;243;207m█[0m[38;2;254;244;211m█[0m[38;2;121;103;91m█[0m[38;2;75;57;54m█[0m[38;2;228;225;224m█[0m[38;2;246;245;247m█[0m[38;2;229;225;225m█[0m[38;2;98;80;79m█[0m[38;2;48;27;22m█[0m[38;2;185;171;147m█[0m[38;2;255;247;215m█[0m[38;2;251;240;208m█████████[0m[38;2;251;241;207m█[0m[38;2;254;245;211m█[0m[38;2;203;189;164m█[0m[38;2;118;103;89m█[0m[38;2;163;154;147m█[0m[38;2;177;171;165m█[0m[38;2;153;143;137m█[0m[38;2;119;102;88m█[0m[38;2;204;192;166m█[0m[38;2;254;244;212m█[0m[38;2;251;240;208m█████[0m[38;2;252;241;208m█[0m[38;2;246;234;203m█[0m[38;2;181;169;140m█[0m[38;2;252;241;209m█[0m[38;2;251;240;208m██████████[0m[38;2;255;251;215m█[0m[38;2;186;171;151m█[0m[38;2;110;82;64m█[0m[38;2;238;202;160m█[0m[38;2;249;209;165m█[0m[38;2;246;205;161m█[0m[38;2;246;205;160m█[0m[38;2;247;206;162m█[0m[38;2;247;206;161m█[0m[38;2;246;206;161m█[0m[38;2;246;205;159m█[0m[38;2;247;204;158m█[0m[38;2;247;204;160m█[0m[38;2;245;205;159m█[0m[38;2;245;204;158m█[0m");
	$display("[38;2;245;201;154m█[0m[38;2;246;202;155m█[0m[38;2;247;203;156m█[0m[38;2;246;202;156m█[0m[38;2;246;203;156m█[0m[38;2;246;205;156m█[0m[38;2;247;206;158m█[0m[38;2;247;205;160m█[0m[38;2;247;205;162m█[0m[38;2;247;206;163m█[0m[38;2;247;205;163m█[0m[38;2;248;206;164m█[0m[38;2;250;208;165m█[0m[38;2;229;197;164m█[0m[38;2;161;156;149m█[0m[38;2;235;203;165m█[0m[38;2;104;76;62m█[0m[38;2;136;120;104m█[0m[38;2;255;248;217m█[0m[38;2;251;241;207m█[0m[38;2;251;240;208m████[0m[38;2;251;241;207m█[0m[38;2;251;241;208m█[0m[38;2;251;230;208m█[0m[38;2;251;214;208m█[0m[38;2;245;202;204m█[0m[38;2;245;198;205m█[0m[38;2;248;200;205m█[0m[38;2;244;197;201m█[0m[38;2;244;197;202m█[0m[38;2;243;198;203m█[0m[38;2;244;199;202m█[0m[38;2;245;209;204m█[0m[38;2;248;229;207m█[0m[38;2;253;244;211m█[0m[38;2;122;104;90m█[0m[38;2;53;33;29m█[0m[38;2;107;90;88m█[0m[38;2;113;101;98m█[0m[38;2;96;79;75m█[0m[38;2;55;33;29m█[0m[38;2;55;35;32m█[0m[38;2;192;178;154m█[0m[38;2;255;246;214m█[0m[38;2;251;240;208m█████████[0m[38;2;253;243;210m█[0m[38;2;237;225;194m█[0m[38;2;74;54;47m█[0m[38;2;68;51;50m█[0m[38;2;202;196;197m█[0m[38;2;235;232;234m█[0m[38;2;212;204;207m█[0m[38;2;72;51;50m█[0m[38;2;63;44;35m█[0m[38;2;220;208;180m█[0m[38;2;254;244;212m█[0m[38;2;251;240;208m██[0m[38;2;251;241;208m███[0m[38;2;252;242;208m█[0m[38;2;254;243;211m█[0m[38;2;251;240;208m███████████[0m[38;2;251;241;207m█[0m[38;2;255;249;217m█[0m[38;2;150;134;117m█[0m[38;2;142;111;88m█[0m[38;2;252;213;170m█[0m[38;2;247;206;164m█[0m[38;2;247;205;163m█[0m[38;2;248;206;163m█[0m[38;2;247;206;163m█[0m[38;2;246;205;160m█[0m[38;2;246;204;157m█[0m[38;2;247;204;157m█[0m[38;2;247;205;158m█[0m[38;2;246;204;157m█[0m[38;2;245;203;156m█[0m");
	$display("[38;2;246;202;153m█[0m[38;2;245;201;152m█[0m[38;2;247;203;155m█[0m[38;2;246;204;156m██[0m[38;2;245;204;155m█[0m[38;2;245;205;156m█[0m[38;2;246;204;157m█[0m[38;2;247;206;161m█[0m[38;2;248;206;165m█[0m[38;2;247;206;164m█[0m[38;2;247;205;163m█[0m[38;2;249;208;163m█[0m[38;2;180;166;150m█[0m[38;2;195;179;162m█[0m[38;2;186;151;123m█[0m[38;2;73;50;43m█[0m[38;2;231;219;190m█[0m[38;2;254;245;210m█[0m[38;2;251;241;207m█[0m[38;2;251;240;208m████[0m[38;2;251;239;208m█[0m[38;2;251;217;211m█[0m[38;2;227;180;189m█[0m[38;2;203;155;164m█[0m[38;2;245;196;205m█[0m[38;2;240;192;201m█[0m[38;2;208;164;170m█[0m[38;2;244;196;203m█[0m[38;2;243;195;202m█[0m[38;2;239;191;198m█[0m[38;2;246;197;205m█[0m[38;2;250;199;210m█[0m[38;2;245;196;203m█[0m[38;2;248;219;206m█[0m[38;2;239;229;198m█[0m[38;2;168;155;132m█[0m[38;2;144;129;115m█[0m[38;2;142;128;117m█[0m[38;2;131;116;105m█[0m[38;2;134;117;103m█[0m[38;2;199;186;161m█[0m[38;2;253;243;210m█[0m[38;2;252;241;209m█[0m[38;2;251;240;208m███[0m[38;2;254;243;211m██[0m[38;2;251;240;208m████[0m[38;2;253;242;209m█[0m[38;2;241;230;200m█[0m[38;2;95;78;67m█[0m[38;2;58;39;35m█[0m[38;2;101;85;81m█[0m[38;2;110;94;92m█[0m[38;2;94;76;74m█[0m[38;2;54;32;30m█[0m[38;2;76;58;49m█[0m[38;2;225;215;184m█[0m[38;2;255;246;211m█[0m[38;2;251;241;208m█[0m[38;2;251;238;207m█[0m[38;2;250;236;206m█[0m[38;2;250;234;207m█[0m[38;2;250;233;207m█[0m[38;2;249;234;206m█[0m[38;2;251;237;207m█[0m[38;2;251;240;208m█[0m[38;2;251;242;208m█[0m[38;2;251;241;208m█[0m[38;2;251;240;208m█████████[0m[38;2;253;242;209m█[0m[38;2;244;235;205m█[0m[38;2;107;83;70m█[0m[38;2;209;173;136m█[0m[38;2;250;210;168m█[0m[38;2;247;206;164m█[0m[38;2;246;204;162m█[0m[38;2;246;204;161m█[0m[38;2;245;203;157m█[0m[38;2;245;203;155m█[0m[38;2;247;205;156m██[0m[38;2;245;203;155m█[0m[38;2;245;202;155m█[0m");
	$display("[38;2;246;202;155m█[0m[38;2;245;202;155m█[0m[38;2;246;203;156m█[0m[38;2;246;204;156m█[0m[38;2;247;206;158m█[0m[38;2;246;205;157m█[0m[38;2;246;205;156m█[0m[38;2;246;203;155m█[0m[38;2;246;205;158m█[0m[38;2;247;206;162m█[0m[38;2;248;207;163m█[0m[38;2;249;207;164m█[0m[38;2;235;204;166m█[0m[38;2;155;150;142m█[0m[38;2;227;198;171m█[0m[38;2;103;74;62m█[0m[38;2;129;112;96m█[0m[38;2;255;249;214m█[0m[38;2;251;241;207m██[0m[38;2;251;240;208m███[0m[38;2;252;242;210m█[0m[38;2;249;219;209m█[0m[38;2;193;149;156m█[0m[38;2;174;133;138m█[0m[38;2;232;185;192m█[0m[38;2;220;175;182m█[0m[38;2;160;120;126m█[0m[38;2;214;169;176m█[0m[38;2;224;178;186m█[0m[38;2;167;125;131m█[0m[38;2;227;181;189m█[0m[38;2;249;200;209m█[0m[38;2;194;150;157m█[0m[38;2;231;183;192m█[0m[38;2;246;198;204m█[0m[38;2;251;234;207m█[0m[38;2;255;250;214m█[0m[38;2;253;243;209m█[0m[38;2;247;236;202m█[0m[38;2;249;239;205m█[0m[38;2;255;247;214m█[0m[38;2;255;247;213m█[0m[38;2;249;238;206m█[0m[38;2;249;239;207m█[0m[38;2;252;242;209m█[0m[38;2;251;240;208m█[0m[38;2;253;242;210m█[0m[38;2;229;217;188m█[0m[38;2;231;219;189m█[0m[38;2;252;241;209m█[0m[38;2;251;240;208m██[0m[38;2;251;241;208m█[0m[38;2;255;246;212m█[0m[38;2;254;244;210m█[0m[38;2;235;224;194m█[0m[38;2;164;150;129m█[0m[38;2;142;129;115m█[0m[38;2;143;131;120m█[0m[38;2;126;111;99m█[0m[38;2;139;123;107m█[0m[38;2;223;211;185m█[0m[38;2;254;237;211m█[0m[38;2;252;223;208m█[0m[38;2;246;209;204m█[0m[38;2;246;202;204m█[0m[38;2;248;201;205m█[0m[38;2;249;201;207m█[0m[38;2;245;197;204m█[0m[38;2;245;198;204m█[0m[38;2;249;203;206m█[0m[38;2;246;206;204m█[0m[38;2;247;217;204m█[0m[38;2;250;234;207m█[0m[38;2;252;242;209m█[0m[38;2;251;240;208m█████████[0m[38;2;255;250;215m█[0m[38;2;173;157;140m█[0m[38;2;136;104;82m█[0m[38;2;252;210;164m█[0m[38;2;246;204;159m█[0m[38;2;245;204;158m█[0m[38;2;246;205;159m█[0m[38;2;244;203;157m█[0m[38;2;242;200;154m█[0m[38;2;242;199;153m█[0m[38;2;240;197;151m█[0m[38;2;236;192;146m█[0m[38;2;236;192;145m█[0m");
	$display("[38;2;246;201;151m██[0m[38;2;245;201;153m█[0m[38;2;246;202;155m█[0m[38;2;246;204;157m█[0m[38;2;247;206;160m███[0m[38;2;247;207;161m█[0m[38;2;248;206;160m█[0m[38;2;247;205;159m█[0m[38;2;250;208;161m█[0m[38;2;220;192;163m█[0m[38;2;165;158;148m█[0m[38;2;225;190;158m█[0m[38;2;70;43;37m█[0m[38;2;183;169;144m█[0m[38;2;255;248;214m█[0m[38;2;251;240;208m█████[0m[38;2;252;242;210m█[0m[38;2;243;208;204m█[0m[38;2;210;163;170m█[0m[38;2;248;199;205m█[0m[38;2;225;179;184m█[0m[38;2;147;108;112m█[0m[38;2;231;185;193m█[0m[38;2;230;183;191m█[0m[38;2;144;104;110m█[0m[38;2;226;179;187m█[0m[38;2;253;204;213m█[0m[38;2;177;135;141m█[0m[38;2;154;116;121m█[0m[38;2;244;197;205m█[0m[38;2;244;197;204m█[0m[38;2;248;230;206m█[0m[38;2;252;241;208m█[0m[38;2;251;240;208m█[0m[38;2;252;241;209m██[0m[38;2;251;241;207m█[0m[38;2;254;245;210m█[0m[38;2;211;200;171m█[0m[38;2;143;130;109m█[0m[38;2;242;233;202m█[0m[38;2;255;245;213m█[0m[38;2;249;240;209m█[0m[38;2;107;91;78m█[0m[38;2;118;103;84m█[0m[38;2;255;250;218m█[0m[38;2;255;247;213m█[0m[38;2;255;247;212m█[0m[38;2;253;242;211m█[0m[38;2;200;189;160m█[0m[38;2;246;235;203m█[0m[38;2;254;244;209m█[0m[38;2;255;248;214m█[0m[38;2;253;242;208m█[0m[38;2;246;235;202m█[0m[38;2;249;239;205m█[0m[38;2;255;245;216m█[0m[38;2;253;218;211m█[0m[38;2;239;194;198m█[0m[38;2;191;147;153m█[0m[38;2;217;168;178m█[0m[38;2;253;202;212m█[0m[38;2;226;178;187m█[0m[38;2;177;134;141m█[0m[38;2;233;184;193m█[0m[38;2;250;202;210m█[0m[38;2;217;169;177m█[0m[38;2;236;186;196m█[0m[38;2;248;196;207m█[0m[38;2;249;202;207m█[0m[38;2;247;220;204m█[0m[38;2;251;240;209m█[0m[38;2;251;240;208m████████[0m[38;2;254;244;209m█[0m[38;2;228;217;190m█[0m[38;2;106;78;60m█[0m[38;2;234;192;148m█[0m[38;2;244;201;154m█[0m[38;2;244;202;154m█[0m[38;2;245;203;156m█[0m[38;2;246;205;159m██[0m[38;2;246;204;159m███[0m[38;2;245;202;158m█[0m");
	$display("[38;2;246;201;152m█[0m[38;2;247;202;152m█[0m[38;2;245;201;152m█[0m[38;2;246;203;153m█[0m[38;2;246;204;157m█[0m[38;2;247;206;160m██[0m[38;2;246;205;160m█[0m[38;2;246;204;159m█[0m[38;2;245;203;157m█[0m[38;2;244;202;154m█[0m[38;2;247;205;156m█[0m[38;2;206;181;155m█[0m[38;2;178;165;152m█[0m[38;2;213;177;141m█[0m[38;2;66;41;35m█[0m[38;2;208;194;170m█[0m[38;2;255;246;212m█[0m[38;2;251;240;208m█████[0m[38;2;251;241;208m█[0m[38;2;250;230;208m█[0m[38;2;249;205;206m█[0m[38;2;248;197;204m█[0m[38;2;226;178;184m█[0m[38;2;230;181;190m█[0m[38;2;254;203;213m█[0m[38;2;194;149;156m█[0m[38;2;205;159;167m█[0m[38;2;252;202;211m█[0m[38;2;246;198;206m█[0m[38;2;207;161;169m█[0m[38;2;238;190;199m█[0m[38;2;246;196;206m█[0m[38;2;245;210;205m█[0m[38;2;250;240;208m█[0m[38;2;251;240;208m█████[0m[38;2;252;241;208m█[0m[38;2;249;238;207m█[0m[38;2;192;181;155m█[0m[38;2;163;150;131m█[0m[38;2;123;107;93m█[0m[38;2;91;71;60m█[0m[38;2;61;38;32m█[0m[38;2;69;46;40m█[0m[38;2;143;127;107m█[0m[38;2;200;188;162m█[0m[38;2;204;193;167m█[0m[38;2;160;145;126m█[0m[38;2;129;114;93m█[0m[38;2;246;235;204m█[0m[38;2;252;242;208m█[0m[38;2;251;240;208m██[0m[38;2;252;241;209m█[0m[38;2;252;242;210m█[0m[38;2;249;218;210m█[0m[38;2;233;185;193m█[0m[38;2;160;121;125m█[0m[38;2;205;162;169m█[0m[38;2;248;199;208m█[0m[38;2;205;159;166m█[0m[38;2;147;106;112m█[0m[38;2;221;175;183m█[0m[38;2;247;198;207m█[0m[38;2;176;133;140m█[0m[38;2;172;130;136m█[0m[38;2;243;193;202m█[0m[38;2;242;194;202m█[0m[38;2;179;136;142m█[0m[38;2;232;184;190m█[0m[38;2;249;227;207m█[0m[38;2;251;243;207m█[0m[38;2;251;240;208m███████[0m[38;2;252;241;207m█[0m[38;2;250;239;208m█[0m[38;2;109;88;72m█[0m[38;2;209;172;134m█[0m[38;2;243;201;157m█[0m[38;2;237;196;152m█[0m[38;2;239;197;152m█[0m[38;2;241;198;153m█[0m[38;2;244;201;156m█[0m[38;2;246;205;159m██[0m[38;2;246;205;157m█[0m[38;2;246;204;157m█[0m");
	$display("[38;2;247;203;155m█[0m[38;2;246;202;155m█[0m[38;2;246;203;156m█[0m[38;2;246;203;157m█[0m[38;2;244;202;155m█[0m[38;2;242;201;153m█[0m[38;2;242;201;154m█[0m[38;2;242;201;155m███[0m[38;2;244;202;157m█[0m[38;2;248;205;158m█[0m[38;2;207;185;157m█[0m[38;2;185;170;152m█[0m[38;2;218;178;141m█[0m[38;2;67;41;36m█[0m[38;2;210;195;173m█[0m[38;2;255;246;212m█[0m[38;2;251;240;208m█████[0m[38;2;251;240;207m█[0m[38;2;251;242;207m█[0m[38;2;251;236;209m█[0m[38;2;248;220;205m█[0m[38;2;248;208;205m█[0m[38;2;248;202;206m█[0m[38;2;245;197;203m█[0m[38;2;245;196;203m█[0m[38;2;246;197;204m█[0m[38;2;245;196;202m█[0m[38;2;245;198;203m█[0m[38;2;249;206;208m█[0m[38;2;248;210;206m█[0m[38;2;249;224;206m█[0m[38;2;251;239;208m█[0m[38;2;251;241;207m█[0m[38;2;251;240;208m███████[0m[38;2;255;248;214m█[0m[38;2;243;231;203m█[0m[38;2;86;61;54m█[0m[38;2;108;70;72m█[0m[38;2;110;74;73m█[0m[38;2;71;42;40m█[0m[38;2;93;58;59m█[0m[38;2;79;51;49m█[0m[38;2;78;54;47m█[0m[38;2;210;197;171m█[0m[38;2;252;241;209m██[0m[38;2;251;240;207m█[0m[38;2;251;240;208m███[0m[38;2;252;242;209m█[0m[38;2;250;221;208m█[0m[38;2;224;176;184m█[0m[38;2;220;173;180m█[0m[38;2;252;201;211m█[0m[38;2;244;196;204m█[0m[38;2;166;124;130m█[0m[38;2;231;183;191m█[0m[38;2;255;205;214m█[0m[38;2;196;151;158m█[0m[38;2;160;119;125m█[0m[38;2;249;202;210m█[0m[38;2;250;201;210m█[0m[38;2;172;129;136m█[0m[38;2;182;138;144m█[0m[38;2;246;198;202m█[0m[38;2;248;225;205m█[0m[38;2;252;242;208m█[0m[38;2;250;241;207m█[0m[38;2;251;240;208m██████[0m[38;2;251;241;207m█[0m[38;2;254;243;213m█[0m[38;2;117;96;82m█[0m[38;2;205;166;133m█[0m[38;2;252;211;164m█[0m[38;2;246;205;159m█[0m[38;2;246;204;159m█[0m[38;2;246;203;158m█[0m[38;2;245;205;159m█[0m[38;2;246;206;160m█[0m[38;2;246;204;158m█[0m[38;2;246;203;157m██[0m");
	$display("[38;2;246;203;155m█[0m[38;2;245;202;153m█[0m[38;2;246;202;155m█[0m[38;2;245;202;156m█[0m[38;2;244;201;154m█[0m[38;2;245;202;154m█[0m[38;2;246;202;155m█[0m[38;2;246;203;156m█[0m[38;2;246;204;157m█[0m[38;2;245;205;157m█[0m[38;2;244;204;156m█[0m[38;2;247;205;156m█[0m[38;2;217;191;158m█[0m[38;2;171;159;147m█[0m[38;2;228;189;151m█[0m[38;2;74;47;39m█[0m[38;2;192;177;155m█[0m[38;2;255;247;214m█[0m[38;2;251;240;208m███████[0m[38;2;251;241;207m█[0m[38;2;251;242;208m█[0m[38;2;251;240;208m█[0m[38;2;251;237;209m█[0m[38;2;250;232;208m█[0m[38;2;250;230;207m█[0m[38;2;250;229;207m█[0m[38;2;250;230;207m█[0m[38;2;251;234;208m█[0m[38;2;251;239;209m█[0m[38;2;251;241;208m█[0m[38;2;252;242;208m█[0m[38;2;251;240;208m█████████[0m[38;2;254;244;211m█[0m[38;2;223;211;183m█[0m[38;2;112;75;73m█[0m[38;2;230;167;181m█[0m[38;2;214;154;168m█[0m[38;2;184;129;142m█[0m[38;2;232;168;184m█[0m[38;2;169;120;128m█[0m[38;2;96;77;67m█[0m[38;2;253;243;210m█[0m[38;2;252;243;209m█[0m[38;2;251;240;208m███████[0m[38;2;251;219;208m█[0m[38;2;248;201;207m█[0m[38;2;245;195;204m█[0m[38;2;245;194;204m█[0m[38;2;245;195;205m█[0m[38;2;247;196;207m█[0m[38;2;247;195;206m█[0m[38;2;231;181;191m█[0m[38;2;240;190;199m█[0m[38;2;247;196;206m█[0m[38;2;245;195;204m█[0m[38;2;229;182;189m█[0m[38;2;248;203;207m█[0m[38;2;248;221;206m█[0m[38;2;251;240;208m█████████[0m[38;2;251;241;207m█[0m[38;2;254;244;213m█[0m[38;2;116;95;81m█[0m[38;2;202;162;128m█[0m[38;2;251;210;162m█[0m[38;2;246;204;159m█[0m[38;2;246;205;159m█[0m[38;2;247;205;159m█[0m[38;2;246;205;158m█[0m[38;2;247;204;157m█[0m[38;2;247;203;157m██[0m[38;2;246;202;156m█[0m");
	$display("[38;2;244;202;153m█[0m[38;2;245;201;152m█[0m[38;2;246;202;154m█[0m[38;2;246;202;155m█████[0m[38;2;246;203;155m█[0m[38;2;246;204;156m██[0m[38;2;248;205;157m█[0m[38;2;229;196;159m█[0m[38;2;153;149;141m█[0m[38;2;230;196;159m█[0m[38;2;96;67;54m█[0m[38;2;150;135;115m█[0m[38;2;255;249;215m█[0m[38;2;251;240;208m██████████[0m[38;2;251;241;208m███████[0m[38;2;251;240;208m██████████[0m[38;2;251;240;207m█[0m[38;2;255;245;211m█[0m[38;2;222;210;181m█[0m[38;2;84;52;48m█[0m[38;2;200;142;154m█[0m[38;2;232;165;183m█[0m[38;2;237;168;187m█[0m[38;2;216;153;170m█[0m[38;2;102;66;70m█[0m[38;2;163;148;129m█[0m[38;2;255;247;214m█[0m[38;2;251;240;208m███████[0m[38;2;251;241;207m█[0m[38;2;252;242;208m█[0m[38;2;251;236;208m█[0m[38;2;249;226;207m█[0m[38;2;248;219;208m█[0m[38;2;248;216;206m█[0m[38;2;247;213;205m█[0m[38;2;247;212;205m█[0m[38;2;249;214;206m█[0m[38;2;249;216;205m█[0m[38;2;248;218;206m█[0m[38;2;248;223;207m█[0m[38;2;251;232;209m█[0m[38;2;251;238;208m█[0m[38;2;252;242;208m█[0m[38;2;251;240;208m█████████[0m[38;2;252;242;208m█[0m[38;2;247;237;207m█[0m[38;2;100;77;63m█[0m[38;2;205;164;128m█[0m[38;2;249;207;158m█[0m[38;2;246;202;156m█[0m[38;2;247;203;157m█[0m[38;2;246;203;157m█[0m[38;2;246;202;155m██[0m[38;2;247;203;156m█[0m[38;2;246;202;155m██[0m");
	$display("[38;2;244;199;150m█[0m[38;2;244;200;152m██[0m[38;2;245;201;153m█[0m[38;2;245;201;154m█[0m[38;2;246;202;155m████[0m[38;2;245;203;155m█[0m[38;2;245;202;155m█[0m[38;2;246;203;154m█[0m[38;2;242;204;162m█[0m[38;2;153;151;149m█[0m[38;2;207;184;159m█[0m[38;2;151;117;95m█[0m[38;2;93;73;59m█[0m[38;2;250;240;207m█[0m[38;2;252;241;209m█[0m[38;2;251;240;208m███████████████████████████[0m[38;2;253;244;211m█[0m[38;2;159;146;121m█[0m[38;2;144;128;110m█[0m[38;2;134;107;99m█[0m[38;2;143;108;105m█[0m[38;2;147;111;108m█[0m[38;2;134;105;98m█[0m[38;2;176;163;142m█[0m[38;2;250;240;208m█[0m[38;2;252;241;208m█[0m[38;2;251;240;208m█████████[0m[38;2;251;241;208m██[0m[38;2;251;242;208m███[0m[38;2;251;242;207m█[0m[38;2;251;242;208m████[0m[38;2;251;241;208m█[0m[38;2;251;240;208m███████████[0m[38;2;254;246;211m█[0m[38;2;217;205;178m█[0m[38;2;77;51;39m█[0m[38;2;222;179;141m█[0m[38;2;247;205;155m█[0m[38;2;245;201;151m█[0m[38;2;246;202;153m█[0m[38;2;246;202;154m█[0m[38;2;246;202;153m█[0m[38;2;246;202;154m██[0m[38;2;245;201;154m█[0m[38;2;244;200;152m█[0m");
	$display("[38;2;245;200;152m█[0m[38;2;245;202;153m█[0m[38;2;245;201;151m█[0m[38;2;245;202;152m█[0m[38;2;246;202;154m█[0m[38;2;245;201;154m██[0m[38;2;246;202;155m██[0m[38;2;247;203;156m█[0m[38;2;246;202;155m█[0m[38;2;246;204;156m█[0m[38;2;251;210;161m█[0m[38;2;184;172;157m█[0m[38;2;162;155;150m█[0m[38;2;204;169;134m█[0m[38;2;68;41;34m█[0m[38;2;196;183;158m█[0m[38;2;255;248;215m█[0m[38;2;251;240;208m██████████████████████████[0m[38;2;251;241;208m█[0m[38;2;252;243;210m█[0m[38;2;139;125;104m█[0m[38;2;208;196;171m█[0m[38;2;251;242;213m█[0m[38;2;235;226;194m█[0m[38;2;231;222;189m█[0m[38;2;246;237;204m█[0m[38;2;255;248;214m█[0m[38;2;252;241;208m█[0m[38;2;251;240;208m████████████████████████████████[0m[38;2;255;250;215m█[0m[38;2;153;138;120m█[0m[38;2;86;56;42m█[0m[38;2;240;198;151m█[0m[38;2;246;204;155m█[0m[38;2;245;201;152m█[0m[38;2;246;201;151m█[0m[38;2;245;201;152m███[0m[38;2;244;201;152m█[0m[38;2;245;201;152m██[0m");
	$display("[38;2;245;202;152m█[0m[38;2;246;203;153m█[0m[38;2;246;202;152m█[0m[38;2;246;201;152m█[0m[38;2;246;201;153m█[0m[38;2;245;201;154m██[0m[38;2;245;203;155m█[0m[38;2;246;204;156m█[0m[38;2;248;204;157m█[0m[38;2;246;203;157m█[0m[38;2;239;196;154m█[0m[38;2;231;187;143m█[0m[38;2;208;176;145m█[0m[38;2;140;140;143m█[0m[38;2;198;176;151m█[0m[38;2;131;100;84m█[0m[38;2;91;73;62m█[0m[38;2;245;234;202m█[0m[38;2;253;243;209m█[0m[38;2;251;240;208m██████████████████████████[0m[38;2;252;241;209m█[0m[38;2;244;233;202m█[0m[38;2;193;181;155m█[0m[38;2;206;194;168m█[0m[38;2;244;234;203m█[0m[38;2;254;245;210m█[0m[38;2;252;241;208m█[0m[38;2;251;240;208m█████████████████████████████████[0m[38;2;253;243;211m█[0m[38;2;238;227;195m█[0m[38;2;74;55;48m█[0m[38;2;139;106;79m█[0m[38;2;246;202;153m█[0m[38;2;240;196;147m█[0m[38;2;242;197;148m█[0m[38;2;244;199;150m█[0m[38;2;245;201;152m█[0m[38;2;246;202;153m█[0m[38;2;246;202;152m██[0m[38;2;248;202;152m██[0m");
	$display("[38;2;247;202;152m█[0m[38;2;246;202;153m█[0m[38;2;246;202;152m█[0m[38;2;246;202;153m█[0m[38;2;246;201;152m█[0m[38;2;246;202;153m█[0m[38;2;248;203;152m█[0m[38;2;246;200;149m█[0m[38;2;237;192;145m█[0m[38;2;221;179;135m█[0m[38;2;211;169;128m█[0m[38;2;218;175;136m█[0m[38;2;231;187;146m█[0m[38;2;245;201;155m█[0m[38;2;206;178;152m█[0m[38;2;153;147;140m█[0m[38;2;207;174;141m█[0m[38;2;76;49;39m█[0m[38;2;140;125;106m█[0m[38;2;255;249;216m█[0m[38;2;252;241;209m█[0m[38;2;251;240;208m██████████████████████████[0m[38;2;252;241;209m█[0m[38;2;255;245;213m█[0m[38;2;251;240;208m█[0m[38;2;250;239;207m█[0m[38;2;251;240;208m███████████████████████████████████[0m[38;2;255;248;215m█[0m[38;2;144;128;111m█[0m[38;2;62;39;30m█[0m[38;2;214;175;135m█[0m[38;2;247;200;149m█[0m[38;2;243;197;149m█[0m[38;2;242;199;149m█[0m[38;2;242;198;149m█[0m[38;2;242;196;147m█[0m[38;2;243;197;148m█[0m[38;2;244;197;148m█[0m[38;2;244;198;149m█[0m[38;2;245;199;150m█[0m[38;2;246;200;150m█[0m");
	$display("[38;2;247;202;153m█[0m[38;2;245;202;153m█[0m[38;2;247;203;155m█[0m[38;2;247;203;156m█[0m[38;2;246;202;155m█[0m[38;2;239;194;150m█[0m[38;2;225;180;137m█[0m[38;2;213;167;124m█[0m[38;2;215;170;128m█[0m[38;2;227;185;139m█[0m[38;2;242;198;152m█[0m[38;2;248;206;159m█[0m[38;2;248;206;158m█[0m[38;2;243;201;153m█[0m[38;2;242;198;150m█[0m[38;2;194;171;144m█[0m[38;2;175;160;146m█[0m[38;2;183;153;124m█[0m[38;2;70;47;34m█[0m[38;2;162;147;128m█[0m[38;2;255;248;214m█[0m[38;2;253;244;209m█[0m[38;2;251;240;208m███████████████████████████████████████████████████████████████[0m[38;2;255;250;216m█[0m[38;2;189;175;151m█[0m[38;2;57;35;27m█[0m[38;2;161;126;98m█[0m[38;2;249;207;157m█[0m[38;2;244;200;151m█[0m[38;2;244;198;149m█[0m[38;2;241;196;147m█[0m[38;2;241;195;146m█[0m[38;2;243;197;147m█[0m[38;2;246;199;150m█[0m[38;2;244;196;147m█[0m[38;2;242;195;146m█[0m[38;2;242;194;145m█[0m[38;2;242;195;146m█[0m");
	$display("[38;2;246;200;151m█[0m[38;2;244;199;150m█[0m[38;2;239;195;146m█[0m[38;2;231;186;141m█[0m[38;2;224;179;138m█[0m[38;2;226;181;140m█[0m[38;2;232;188;144m█[0m[38;2;240;194;145m█[0m[38;2;246;198;148m█[0m[38;2;247;200;150m█[0m[38;2;246;200;151m█[0m[38;2;243;198;152m█[0m[38;2;240;197;149m█[0m[38;2;236;193;145m█[0m[38;2;235;192;144m█[0m[38;2;242;197;148m█[0m[38;2;221;186;149m█[0m[38;2;201;179;149m█[0m[38;2;177;146;120m█[0m[38;2;69;46;36m█[0m[38;2;136;121;104m█[0m[38;2;243;235;201m█[0m[38;2;255;248;215m█[0m[38;2;252;241;209m█[0m[38;2;251;240;208m███████████████████████████████████████████████████████████[0m[38;2;252;242;208m█[0m[38;2;255;250;216m█[0m[38;2;194;182;159m█[0m[38;2;65;43;35m█[0m[38;2;141;108;83m█[0m[38;2;248;205;158m█[0m[38;2;247;203;155m█[0m[38;2;245;202;154m█[0m[38;2;245;201;152m█[0m[38;2;244;198;149m█[0m[38;2;242;196;147m█[0m[38;2;241;195;146m██[0m[38;2;242;194;145m██[0m[38;2;245;197;148m█[0m[38;2;246;198;149m█[0m");
	$display("[38;2;234;189;140m█[0m[38;2;232;188;139m█[0m[38;2;233;189;140m█[0m[38;2;237;194;145m█[0m[38;2;244;200;153m█[0m[38;2;247;203;154m█[0m[38;2;245;202;152m█[0m[38;2;245;199;150m█[0m[38;2;243;196;147m█[0m[38;2;240;194;145m█[0m[38;2;239;193;144m█[0m[38;2;239;194;146m█[0m[38;2;238;194;146m█[0m[38;2;239;194;147m█[0m[38;2;241;196;149m█[0m[38;2;242;196;148m█[0m[38;2;240;194;145m█[0m[38;2;230;189;140m█[0m[38;2;233;192;148m█[0m[38;2;208;165;125m█[0m[38;2;102;71;57m█[0m[38;2;89;71;57m█[0m[38;2;190;178;152m█[0m[38;2;249;239;207m█[0m[38;2;255;246;212m█[0m[38;2;251;241;208m█[0m[38;2;251;240;208m████████████████████████████████████████████████████████[0m[38;2;254;244;211m█[0m[38;2;250;241;210m█[0m[38;2;165;151;133m█[0m[38;2;75;51;42m█[0m[38;2;150;115;88m█[0m[38;2;237;195;149m█[0m[38;2;244;201;154m█[0m[38;2;246;202;154m█[0m[38;2;245;201;153m█[0m[38;2;246;200;152m█[0m[38;2;246;200;151m█[0m[38;2;246;199;151m██[0m[38;2;245;198;149m█[0m[38;2;244;196;147m█[0m[38;2;242;194;145m█[0m[38;2;244;196;148m██[0m");
	$display("[38;2;241;194;146m█[0m[38;2;244;197;148m█[0m[38;2;245;200;151m█[0m[38;2;246;201;152m█[0m[38;2;245;200;150m█[0m[38;2;245;199;150m█[0m[38;2;242;196;147m█[0m[38;2;238;192;143m█[0m[38;2;240;193;145m█[0m[38;2;241;195;146m█[0m[38;2;241;196;147m█[0m[38;2;242;196;147m█[0m[38;2;244;198;149m█[0m[38;2;244;197;148m█[0m[38;2;238;192;143m█[0m[38;2;236;191;142m█[0m[38;2;237;192;143m█[0m[38;2;234;188;138m█[0m[38;2;238;191;142m█[0m[38;2;247;201;152m█[0m[38;2;243;201;153m█[0m[38;2;162;126;96m█[0m[38;2;76;49;37m█[0m[38;2;111;93;77m█[0m[38;2;196;183;159m█[0m[38;2;249;239;207m█[0m[38;2;251;241;208m█[0m[38;2;251;240;208m██████████████████████████████████████████████████████[0m[38;2;253;243;210m█[0m[38;2;221;211;183m█[0m[38;2;118;102;89m█[0m[38;2;107;77;59m█[0m[38;2;204;164;126m█[0m[38;2;238;194;147m█[0m[38;2;218;174;128m█[0m[38;2;218;173;129m█[0m[38;2;231;185;137m█[0m[38;2;241;195;146m█[0m[38;2;244;198;149m█[0m[38;2;245;199;150m█[0m[38;2;245;198;149m███[0m[38;2;245;197;148m█[0m[38;2;245;197;149m█[0m[38;2;247;199;151m█[0m[38;2;245;197;149m█[0m");
    $display ("--------------------------------------------------------------------");
    $display ("                         Congratulations!                           ");
    $display ("                  You have passed all patterns!                     ");
    $display ("                  Your execution cycles = %5d cycles                ", total_latency);
	$display ("                  Your clock period = %.1f ns                       ", CYCLE);
    $display ("                  Total Latency = %.1f ns                           ", total_latency*CYCLE);
    $display ("--------------------------------------------------------------------");     
    repeat(2)@(negedge clk);
    $finish;
end endtask

endmodule