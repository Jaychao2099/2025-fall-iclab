//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2025 ICLAB Fall Course
//   Lab09      : RPG
//   Author     : Tzu-Yun Huang
//	 Editor		  : Erh-Yi Tu
//                
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : pseudo_DRAM.sv
//   Module Name : pseudo_DRAM
//   Release version : v2.0 (Release Date: Oct-2025)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`include "Usertype.sv"

module pseudo_DRAM(input clk, INF.DRAM inf);

`protected
):a5QA=&JQD3<+)_c5SbU-5?F0^TWXR<1L[Qf:9>-[5DDJ>DfT^G,):30^F]JWK&
3042D3DKY#MB0R3;])J<;S,a9\7?d.+7?$
`endprotected

//================================================================
// parameters & integer
//================================================================

parameter DRAM_p_r = "../00_TESTBED/DRAM/dram.dat";

parameter DRAM_R_latency = 1;
parameter DRAM_W_latency = 1;
parameter DRAM_B_latency = 1;

`protected
3(FZTVLW<D>=;W9M7-+UGK_f<XS7ObRG9,HfF#6IFaG+>&C&(:GG-)c\D3f#V#HV
97CM<c2B.1eZ=.6G/@(>b)7NPG&S<Q2K0M>C8__=Q:bDg<MM&1CTEAOB5726[]g)
]RLY5UWd,0c1HMI@-6BY4bGJ)^JMb\OT:1H/Z9\T9UD\bY44,Rg&^c@\0?)^R],&
V_(R8],PO/@a=BMV5:IE8fRNZ\-NeJ9#DGafRV\MR8AG+f,B>E(f7,I&>PSUO(TL
HDO/Z(WTdBW-A)3H&IWQU3._+OW_,G9>L1VEFBCG2)C,4PH:WFH(Q.@HK1a<Sc<F
:PE[8LHa8A,c\R<f88_bL.E;#aMB:@+R661QeSQNRDDagfgEOfO=0T-S4f/N6]aO
BWR1TS\e\NAD>cI7^30T+T<b^1C:QB&7035VR;[O9e<WVA>7b9._ObQH2GEGGXP\
5&f2ASUb<[IU7(\RQRa6.@PP8&3@@]>HUad_/^)1Yb#QGC<_7J5/cGKFLNU6I-.#
5PbOM^I7F5Z&R:gg567L3\RN7D02JK[W[<KD#ScU#[(Q:BcIO>=&()e.cR8CL73M
_2JBZEc-fAY=1gHV4_></=Df53a#G64U@4d[TI1MLb&D&WD;Z:g8eN\^cLVE0:?&
Z#H=)a?P:-]e4<URS:4/JX7TU071e[_QT3FPW\O<B(9JU<G.MSD,,4WRJMPLO[V:
B^7:&:UU+b4fS=e#>f&?P,]4We/@+OeZU_f8GIM)MLY]WDWb6W2X/F2aI\#?,X]0
L_>RU?:;:Z/Vb5</R><2e>c_XAX1EWH8M<AH7F/4a6[cRVe__X]bVe.?1fdA&&A2
R]a#Q613X>U:K&Gb/:@EV.,,UBGfWe:?7Kd(M48]:51&dF&MXZ\F&C3RY55\VU&^
gN8[MB=96G=3.[-NP3MJ?KGdPK9)8.b,9@-I42D9LW^J[c1?QAJfON8TQ#+A+YEJ
Q(45Yc9W<+J:VZPKZ[C0O3)),M5S58G</(GB[e_0]R3-JCU&(RbZGV1^Lg]XL.A9
V5e-#7=NU@L+_Q:,4I@U0Y)4;3^JG8K_T=ZPRUS5_V84WI]J/aFB_-TB@(E=;?]G
_U1)RPEN0D2I(8BM_WBEFBd](,d)Pb.W,>Ee+fNC_S]f[bP1_IfZU?f>OJAW[1O7
8BQHKaDC_\7M25>D4;BN8ZRJ]Wdd>dZ<H\[N[9^O&LKFA0MI\A(U)?FSBA&1<]K<
D9/6gD1@FNWP/Q2:XJ9R(_\E.F+#SNZC/O[6L5Y@&@dMeNP(/9\S#f3gM+C:U>^#
a2bN4#gYKV,+3]S>ZS/BC/gEH[LK6(ZY6+IT<MbfM(M[TLTa79MOdg<Fg)W0,RNU
;)7>dULd5a/]eO61LgJ>40d@>M)ea@bCK0.=aPSHbbEFf(.Sb]Q77(<^e3H/T3Sc
>g,^D5TAR8JIU47YW;,[P5AC/3^g8b^-U\=5^.8(Y\9LJL,UKA1AJU\A7d,B/._K
ef:NHJP&N<U:X14Ba0,5]fERAY@aL&c+_C1.;?dX6#Ncd(Va4_./(F3H:-2(&dVP
EHTc2BL2LDJbDZb_\eN(#\9-/Z(.cMe#V,[3/I(]Vb52[,J^165O?(?B\J(K9XS/
[+T:_P9;UCLVPA4a,9V].I(7^b-=X5aZ<<&da:H3_[F=Q1L2WT(^GcR;D_X,>6M7
UA5eH#LQc0F<^Z8;Aa.1;FG3P5(2]Y8=.OUYM+cB+g4WU<6BIU?d[W+79F@=3g\3
L6L=LTg3LK.ff1\-5-J)0J)T9+Y=cJI(b9QEK98)(0:[\2bR7ZQKSSaX/SYSDaD)
YHH]a-+2a3d13IJ)\UQA8(e50b?_d:F9-1I5QPcPB^,F>I#ME3GMd=+FUAZ;5X9)
;7H(+4]^HC6ZG_+C],g354=>RLY.1W+Z=>(R)7S@1\[PR9-bPXU?4Wg2QNcDX,Q6
g+AZ8.3\<U:)+@2+&b5U)fKKA9,Md9KWe;@ZAK1EQ:L],0M9e<Y\a4W]2aP8#8@]
bGK^X=Q0F\5C@Ec:9^[KKQTQ^D?IB<f4E768:3.(L?bg9T(c5;O?CPb@RB&W_+@5
eLM1XYfRdHXY.fF@HFW4,QQ78C.]MOXD\5e\Q44]>>MAU@dR[aBAD,g=OO54<BNI
N?SDV#a(H9Ec:X+\.BaW-&;:)CC</H>gH:)fJP5>R&]Wg2JFeR2B=0H#N_Hd842R
)<:,W/e)[?bQc4N(Y,>X1a4I3Z^,Vdg@+<AKUDd8-de,TUdA3]UgV<\IIY59#HFS
#I6E<KJZ?TDP7)a07OL8@]XV&YK0.fIP9c2KK#J_<N.8bD_3:BeH\4,+2.KN1\+[
O_VG7=SS<],VO&?R>W<]WZ[/YJ@f7C=>^3,E^aF8>4aFFQWa>78J67)7?Hc>P,JT
/6c7Z?:1a#,=<K[9c&18^X0^V-L1_(4V(.RBEUDXS;;+OYXM:1>ROZf4@D)M@[H,
Ag6&MD=W@HcV9PS:e<d8KH@fQd[B?bD=^@UZRL+6M<XMF?,F:=NZEW9\+;4@Eg@X
GS6&Z-DbJZ2XMH4P_d]&W5)d-)/844V^OLR[IMHB1]O3:P,7D3,=ae[V+2]g(^-T
X.QH]g^D@&gWNDE[SJT1b87C0a31SL2T.^fA=5LeGR4.CHI;MKdTXWT?CRQKY5Jb
cbgH9c?fJQQd,BL=-BNWGcG7&1U\-]:L5gI:<\O+G<8KR=a(X/Q@LOOX\9:NX4)e
Q9B5<MfQ/D=\3f4c<+JcX#NY;-@Fg>ZH/G1f@9CY,S6]G\E#]e-,?b.H/MYR.Ra6
]D@CB)a?e&9#VIWLTKO_b-UAE,d/=GH5[Lca^9#;YU20\^TM+&(cU<K1JHQ_dUW1
K?SaE=bB[G@9\6FNI4g-Ra6c1]<(NW4O,R=7E_7<VGHb^#7?0?d73,eV]72&Fc>e
G@X@1)A?+H]Na&&J]TO7;Pg<bMR5SH_,DWgZ^A.L+#dMZ>.d)+gC:V:L[E@9Y9LY
dX:TLF4NI0SMO8f):Y67.V;[NZKMfa=YHE@.QD4f+^cG;@]fC^@R5K[&]].GPQH5
6+]GD2(MA^4(3a<JL:]f+_K5;gG?=)K]VXY/W.,./4?c.J9/L[LfQ?0I_f1GbMH6
^@B96;30N;?=6XR,&bA^6b:\-gHZ#[7<Gb;ZP_EI10RAJX9VLbJGd;6KB=\3@80g
?5&6#MM-aNX[2f#WTSS6b9J.K0:/LgL[5(F[A3#O_SJ:/1&#J(<GN#1_(9][([AN
:J7V7^O)[2)?#X2QY)7Y0E5L#LT.VG=MNW8/#3Y3eC92@XDeJCS\+<042>@IG45N
6D]H^P&>515@fZ#1_4\NVO@3a?ULDOCZXPb7-D(0++f8bU(-Q8Q=<U6NLVL9DGS:
Q]4/72@V7>EG)SVG:1Q+A#T,ZGcaP\)bFC+\)fdd(:9(_8d+RA@YJ;4T4^\/4\ed
BbL2+4>@LB_L@0PWGK[(K7dBV.WEP<R78NI+Z,=W4,Bf^]MFg3E/SL#?ZcU1g0a>
aH&&A?^A7^TM00>LD=TdXY7X?V+aeVVRe<M\b]4JZE29[8^W#AT3#a[78X7J56EV
13P;_e8a:OG.?[JKWCcNaLI(+dFOB)-WBK2V5U?d9V]7V..&6HNb6b[.KD;0[;Y]
e1Z.]3IHg2b#3)c9,=]F_MO&6D^9Wea#0S&6]);>M-Y(>Tf=Bd68X73B12YefaU/
&@Nf\DVg?b-,-(a^Q#^GD<46,/cSQ?^F\M_ZA(6W9+784f-2Pg\-FJ@6T,E#_Q\.
(+B93YH-ZV;/.#,?M@8.J8[=Qdf76_9I0gF.U;4F)[#\TIB8)HL:WXWKS&87LQQ.
8\MF&5+.N.V/RVL0Y.^Q2YV3_^D72H\0IbaG0-aB)UP2@S.@;-.P5J.T3B?@c_.;
^?RV7JR,?6UQ/>/eAb<BW2P,Q[e\&>CB,/46?D@[b1&=a#_U9KBS;4=+_4OOH++1
6KF:@&ed[E-ZT5]T@QC0bZO>+d7K<E1QYVK>WSWMDV(D/GMZ60TS^RKTB[]JFdG6
<g>>G-f99,,X;BD;Z0ZSgZbGBFJ-S=bO0?REOGUd<34=JVW;UT0>cVDCfNE062D1
IaVJc>N<AU@G:X8^QJf60FREB#?6^0>ZTT/Y#@@>Y/)O2?990(]-X]c@AAEGJBG1
(GBKS73<1?]Q1(5KE?g-2)9.GIS;F8C+&a#KV.AX+Ac5Z>CILJWc<fe;/gLN,CT6
(:;(UF4.>9U5\TLOFLO95;4b,3WZ:[([4C:-X-?<Ef;9cD3eY)+dUc4JJ7>QV=3;
+W?b6?E=1E_C6Q]U_IG?D6@BFg>87W(G20O&&RV0>0e[_ET#ELV74G3.>]W9gQ8:
CCP5c#E)62#TEAc7D>;Ob#0B-LJ6EN_C2-;KK1T\NM:JS3a;^0Sf&BAf2/.O9_B4
NeDSXdd[,P\.c]P=D:XL1:B)6G18<:OHA2KH(,MC.If12>-,-AZH7\Ed.D0/#704
\>4;HA1Z>FDNBWQWP)M(gKWR^OXDKcC</B0B:&71D^H68W_B[Na+/CO-8^&d&/3M
Ob@+Z^I#M(RDR?cFCU3V7.C]K#d(D5?d^O<)Ze85]&KYX1cGH[&_B5NT:2YRe5C)
]5?d/A-(XBR^5\4^3B8ON[=e+ML.QIV#4a8V-MFD+dX#J#?Z(R6bGKYZcHAAebSO
6@+(:bH@dX[eS#9;7(0=-/VQ<F0^U5?=S?9OagP2^a2VI^/75UT+1P(;[AJF]X(b
8+&g)bZ^#3IZ?]6X8<#KEK\KTd=YHf\PcRG7;d-gXA706GCY<:VbOKOE=SF<&7fC
E@[(g__#e-b2J[63>HCc>>QXF8Y,UO^^]f5eT65ITP:(MO;..-2U:0:e;&d_f.f3
);/?U=63)348N[(+O5OR8SWf1[4U.HG@=bb;?6]MRR?;4I&=)(ZR\E1D]_;<A>5Z
#8H)WQPC]b7O,_.OY.#]0V:\X1=W>0d,AeO5&G1M>-/OY]17GD9b?3.V3O006QZ9
?>?G.gEOLP9+\,?]&R]#X?(A(@/1(eYb&/U+(@U#^G^b3)9I-L6EI.R?XT]A:PgH
S.UZH[WU#7=9LGRVH6M+<-).Y97U;UL>0>^M(0F\Y6X^K39YZ@Q;/#VI-Zb?H+3b
Fe>7c/c00W=T:ebcQ3Td68b+,L<aN_UJ;;Df:R/W+RW/<U[L6PaG/DJR,W5I/\_1
fD#)^#;H_(2^a@Pecaa(1PfI]08S2\TBd147J&gRQVTP,/_S_:1+BD;fZ;_?+X[(
7>#,4T,#O65C7DED[g)#/WL:3.bea-0/S)ET#\\2TTG2U6DDR22X/fNJEa;E.V_@
<XdN[#SX;/Pd72bfM[LW>FW30=PZWLTH8H@]Z-PK;S2d\,V:XW>;cO#@N,BWY[L\
eNX=C:If,fcMIM@3&)OeAARM-@;8Ra;-7^_VD[A,XFFFTED\8d@SFY19G2KJE=LR
^[KIaAS+7\X)_^cG7I<HP2/C>ZPE+,Cc,[DRC5Wac2Fc(G;I>U]2gZaYgbMR8R)M
TBQQD&UdKZ2ASGM#@5X-ef=<28]-fDb((O6eAJ@CSX]3cQXR2_Qa0?<AW]FJ4=Hc
A<B_GYGc]&N-/7E>CH-4_UM)R_AG10ee^Y:-N^D?,&V,OVH,Ja:OVVI\UU52&K=1
<=RcFY[79Ze-0$
`endprotected
endmodule
