//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2025 ICLAB FALL Course
//   Lab02       : Testbench and Pattern
//   Author      : Ying-Yu (Inyi) Wang
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : v1.0
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`ifdef RTL
    `define CYCLE_TIME 10.0
`endif

`ifdef GATE
    `define CYCLE_TIME 10.0
`endif


module PATTERN(
    // Output signals
	clk,
    rst_n,
	in_valid,
	in,
    // Input signals
    out_valid,
    out
);

//================================================================ 
//   INPUT AND OUTPUT DECLARATION
//================================================================
output reg clk, rst_n, in_valid;
output reg [3:0] in;
input out_valid;
input [3:0] out;

//================================================================
// parameters & integer
//================================================================
real CYCLE = `CYCLE_TIME;
parameter PATNUM = 100;  
integer patcount, total_latency, wait_val_time;
integer i, x, y;
integer in_read, in_hold, out_read, out_hold;

//================================================================
// wire & registers 
//================================================================
reg [6:0] ans, solution;

//================================================================
// clock
//================================================================
initial 
begin
	clk = 0;
end
always #(CYCLE/2.0) clk = ~clk;

//================================================================
// initial
//================================================================
initial 
begin
	//+++++++++++++++++++++++++++++++++++++++++++++++++++
	in_read=$fopen("../00_TESTBED/input.txt","r");
  	out_read=$fopen("../00_TESTBED/output.txt","r");

    // in_read=$fopen("../00_TESTBED/input_1000.txt","r");
  	// out_read=$fopen("../00_TESTBED/output_1000.txt","r");

    // in_read=$fopen("../00_TESTBED/puzzles.txt","r");
  	// out_read=$fopen("../00_TESTBED/solutions.txt","r");

    // in_read=$fopen("../00_TESTBED/input1.txt","r");
  	// out_read=$fopen("../00_TESTBED/output1.txt","r");

    // in_read=$fopen("../00_TESTBED/input_3.txt","r");
  	// out_read=$fopen("../00_TESTBED/output_3.txt","r");
	//+++++++++++++++++++++++++++++++++++++++++++++++++++

	rst_n = 1'b1;
	in_valid = 1'b0;
	in = 'bx;
	force clk = 0;
 	total_latency = 0;
 	
	reset_signal_task;
	
	for(patcount = 1; patcount <= PATNUM; patcount = patcount + 1) 
	begin

        x = 0;
        solution = 'd81;

		input_task;
		wait_out_valid;
		check_ans;
	end	
  	YOU_PASS_task;
end 

always begin	
	if(out_valid===0&&out!=='b0)begin
        $display ("---------------------------------------------------------------------------------------------");
        $display ("             Fail! The out_data should be reset after your out_valid is pulled down.                   ");
        $display ("---------------------------------------------------------------------------------------------");
        repeat(2) #CYCLE;
        $finish;
    end
	else @(negedge clk);
end

// I/O_valid overlap
// always begin	
// 	if(out_valid===1&&in_valid===1)begin
//         $display ("---------------------------------------------------------------------------------------------");
//         $display ("             Fail! The out_valid should not be high when in_valid is high.                    ");
//         $display ("---------------------------------------------------------------------------------------------");
//         $finish;
// 	end
// 	else @(negedge clk);
// end

//================================================================
// task
//================================================================
task reset_signal_task; 
begin 
    #(10);  rst_n=0;
    #(5);
    if((out_valid !== 0)||(out !== 'b0)) 
    begin
        $display ("---------------------------------------------------------------------------------------------");
        $display ("             Fail! Output signals should be 0 after reset at %4t.", $time);
        $display ("---------------------------------------------------------------------------------------------");
        $finish;
    end
      
    #(50);  rst_n=1;
    #(3);  release clk;
end 
endtask

task input_task; 
begin
	// Inputs start from second negtive edge after the begining of clock
    if(patcount=='d1) repeat(2)@(negedge clk);

	// set in_valid and in
    in_valid = 1'b1;
    wait_val_time = 0;
    for(i=0; i<81; i=i+1)
    begin
        in_hold=$fscanf(in_read,"%d",in);
        if (out_valid !== 1) begin
            wait_val_time = wait_val_time + 1;
        end
        @(negedge clk);
    end
    
	// Disable input
    in_valid = 'b0;
    in = 'bx;        
end
endtask

task wait_out_valid; 
begin
    // wait_val_time = 0;
    while(out_valid !== 1) begin
	    wait_val_time = wait_val_time + 1;
	    if(wait_val_time > 1000)
        // if(wait_val_time > 100000)
	    begin
		    $display ("---------------------------------------------------------------------------------------------");
		    $display ("             Fail! The execution latency is over 1000 cycles.");
            // $display ("             Fail! The execution latency is over 100000 cycles.");
		    $display ("---------------------------------------------------------------------------------------------");
		    repeat(2)@(negedge clk);
		    $finish;
	    end
	    @(negedge clk);
    end
    total_latency = total_latency + wait_val_time;
end endtask

task check_ans; 
begin
    // Check the answer here
    
    while(out_valid)
	begin
		
		// out_hold=$fscanf(out_read, "%d", ans);

		if(x>=solution)//x>max-1
		begin
            $display ("---------------------------------------------------------------------------------------------");
            $display ("             Fail! OUT_VALID is over %d cycle(s)", solution);
            $display ("---------------------------------------------------------------------------------------------");
            repeat(9) @(negedge clk);
            $finish;
		end	        
		// if(out!==ans)//complete the if statement here(one statement)
		// begin     
        //     $display ("---------------------------------------------------------------------------------------------");
        //     $display ("             Fail! ANWSER IS WRONG!          ");
        //     $display ("             PATTERN NO.%4d . %4d ",patcount, x+1);
        //     $display ("             Ans:%d  ", ans);//show ans
        //     $display ("             Your output : %d  at %8t ",out, $time);//show output
        //     $display ("---------------------------------------------------------------------------------------------");
        //     repeat(9) @(negedge clk);
        //     $finish;
		// end
		@(negedge clk);	
		// x=x+1;
	end
	
	if(x<solution) 
	begin
		$display ("---------------------------------------------------------------------------------------------");
		$display ("                   Fail! OUT_VALID is less than %d cycle(s)", solution);
		$display ("---------------------------------------------------------------------------------------------");
		repeat(3) @(negedge clk);
		$finish;
	end	
  //+++++++++++++++++++++++++++++++++++++++++++++++
    $display("\033[0;34mPASS PATTERN NO.%4d,\033[m \033[0;32mexecution cycle : %3d\033[m", patcount, wait_val_time);
    repeat(3)@(negedge clk);
end 
endtask

task YOU_PASS_task; 
begin
	display_pass;
    $display ("--------------------------------------------------------------------------------------------------");        
    $display ("                                          Congratulations!!!                         ");
    $display ("                                   You have passed all patterns!                     ");
    $display ("                                   Total lentency : %d cycles                     ", total_latency);
    $display ("--------------------------------------------------------------------------------------------------"); 
	          
         
    #(500);
    $finish;
end
endtask

//Check Ans
always @(posedge clk) begin
    if (out_valid) begin
        out_hold=$fscanf(out_read, "%d", ans);

        if(out!==ans) begin//complete the if statement here(one statement)
            $display ("             \033[0;31mFAIL Pattern NO. %d\033[m         ", patcount);
            display_fail;
            $display ("--------------------------------------------------------------------------------------------------"); 
            $display ("                                Fail! ANWSER IS WRONG!          ");
            $display ("                                PATTERN NO.%4d . %4d ",patcount, x+1);
            $display ("                                Ans:%d  ", ans);//show ans
            $display ("                                Your output : %d  at %8t ",out, $time);//show output
            $display ("--------------------------------------------------------------------------------------------------"); 
            repeat(9) 
            @(negedge clk);
            $finish;
		end
        
        x = x + 1;
        @(negedge clk);
        
    end

end

task display_fail; begin

$display("[38;2;0;0;0m████████████████████████████████████████████████████[0m[38;2;167;163;164m█[0m[38;2;36;34;35m█[0m[38;2;0;0;0m██████████████████████████████████████████████[0m");
$display("[38;2;0;0;0m███████████████████████████████████████████████████[0m[38;2;23;23;23m█[0m[38;2;237;233;221m█[0m[38;2;236;234;222m█[0m[38;2;236;236;224m█[0m[38;2;239;239;229m█[0m[38;2;232;232;222m█[0m[38;2;0;0;0m███████████████████████████████████[0m[38;2;148;148;140m█[0m[38;2;204;200;188m█[0m[38;2;146;145;140m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m██████████████████████████████████████████████████[0m[38;2;0;1;3m█[0m[38;2;199;168;150m█[0m[38;2;213;185;164m█[0m[38;2;220;193;166m█[0m[38;2;221;190;162m█[0m[38;2;222;194;170m█[0m[38;2;217;196;169m█[0m[38;2;204;188;172m█[0m[38;2;218;208;199m█[0m[38;2;0;0;0m████████████████████████████[0m[38;2;0;0;2m█[0m[38;2;51;50;45m█[0m[38;2;241;241;215m█[0m[38;2;238;242;219m█[0m[38;2;242;239;222m█[0m[38;2;244;238;222m█[0m[38;2;241;235;221m█[0m[38;2;233;227;213m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m██████████████████████████████████████████████████[0m[38;2;1;1;3m█[0m[38;2;136;103;70m█[0m[38;2;170;138;100m█[0m[38;2;200;166;139m█[0m[38;2;196;169;140m█[0m[38;2;197;171;148m█[0m[38;2;199;177;156m█[0m[38;2;199;183;158m█[0m[38;2;197;183;170m█[0m[38;2;200;187;181m█[0m[38;2;93;89;88m█[0m[38;2;0;0;0m█████████████████████████[0m[38;2;90;85;79m█[0m[38;2;242;228;215m█[0m[38;2;240;231;214m█[0m[38;2;238;236;215m█[0m[38;2;237;237;211m█[0m[38;2;240;236;209m█[0m[38;2;236;232;205m█[0m[38;2;237;231;209m█[0m[38;2;235;227;208m█[0m[38;2;43;44;38m█[0m[38;2;0;0;2m█[0m[38;2;0;0;0m███[0m");
$display("[38;2;0;0;0m██████████████████████████████████████████████████[0m[38;2;21;16;13m█[0m[38;2;122;96;73m█[0m[38;2;177;150;120m█[0m[38;2;202;174;153m█[0m[38;2;196;174;151m█[0m[38;2;197;176;157m█[0m[38;2;197;180;164m█[0m[38;2;200;173;162m█[0m[38;2;193;171;157m█[0m[38;2;188;172;157m█[0m[38;2;187;173;164m█[0m[38;2;191;184;178m█[0m[38;2;0;0;0m███████████████████████[0m[38;2;92;82;72m█[0m[38;2;186;161;131m█[0m[38;2;224;193;164m█[0m[38;2;241;226;203m█[0m[38;2;241;229;203m█[0m[38;2;235;229;197m█[0m[38;2;240;229;199m██[0m[38;2;237;226;196m█[0m[38;2;229;216;184m█[0m[38;2;222;206;180m█[0m[38;2;1;0;5m█[0m[38;2;0;0;0m███[0m");
$display("[38;2;0;0;0m██████████████████████████████████████████████████[0m[38;2;24;15;8m█[0m[38;2;110;76;39m█[0m[38;2;180;146;119m█[0m[38;2;198;169;153m█[0m[38;2;196;170;155m█[0m[38;2;194;172;159m█[0m[38;2;190;172;162m█[0m[38;2;188;171;163m█[0m[38;2;195;178;170m█[0m[38;2;203;186;178m█[0m[38;2;193;176;166m█[0m[38;2;176;162;153m█[0m[38;2;180;166;157m█[0m[38;2;72;64;62m█[0m[38;2;1;0;2m█[0m[38;2;0;0;0m█████████████████[0m[38;2;0;1;0m█[0m[38;2;2;2;0m█[0m[38;2;114;96;60m█[0m[38;2;166;140;113m█[0m[38;2;225;199;174m█[0m[38;2;229;206;165m█[0m[38;2;237;214;180m█[0m[38;2;235;220;179m█[0m[38;2;233;222;177m█[0m[38;2;240;221;189m██[0m[38;2;235;216;184m█[0m[38;2;225;209;183m█[0m[38;2;202;195;169m█[0m[38;2;93;86;76m█[0m[38;2;0;0;0m███[0m");
$display("[38;2;0;0;0m████████████[0m[38;2;246;4;0m█[0m[38;2;254;1;0m█[0m[38;2;0;5;4m█[0m[38;2;0;0;0m███[0m[38;2;13;0;0m█[0m[38;2;254;1;0m█[0m[38;2;253;1;0m█[0m[38;2;0;0;0m█[0m[38;2;0;2;2m█[0m[38;2;254;1;0m██[0m[38;2;251;2;0m█[0m[38;2;43;0;0m█[0m[38;2;0;0;0m███[0m[38;2;254;2;0m█[0m[38;2;254;1;0m██[0m[38;2;35;0;0m█[0m[38;2;0;0;0m████████████████[0m[38;2;26;19;13m█[0m[38;2;115;74;56m█[0m[38;2;158;122;96m█[0m[38;2;186;155;135m█[0m[38;2;183;165;151m█[0m[38;2;194;176;166m█[0m[38;2;200;181;175m█[0m[38;2;203;186;178m█[0m[38;2;205;188;178m█[0m[38;2;199;183;168m█[0m[38;2;191;174;158m█[0m[38;2;176;162;149m█[0m[38;2;205;190;183m█[0m[38;2;210;199;193m█[0m[38;2;222;215;207m█[0m[38;2;41;40;38m█[0m[38;2;1;0;0m█[0m[38;2;44;43;41m█[0m[38;2;173;168;165m█[0m[38;2;29;28;26m█[0m[38;2;16;15;13m█[0m[38;2;43;43;43m█[0m[38;2;0;0;0m█[0m[38;2;0;0;2m█[0m[38;2;71;72;67m█[0m[38;2;0;0;0m███████[0m[38;2;117;100;70m█[0m[38;2;139;114;84m█[0m[38;2;206;175;155m█[0m[38;2;197;170;140m█[0m[38;2;209;178;147m█[0m[38;2;224;190;153m█[0m[38;2;236;201;163m█[0m[38;2;239;207;168m█[0m[38;2;242;214;175m█[0m[38;2;234;212;171m█[0m[38;2;235;207;168m█[0m[38;2;225;195;159m█[0m[38;2;211;195;162m█[0m[38;2;183;166;138m█[0m[38;2;0;0;2m█[0m[38;2;0;0;0m███[0m");
$display("[38;2;0;0;0m████████████[0m[38;2;251;1;3m█[0m[38;2;254;0;0m█[0m[38;2;0;1;5m█[0m[38;2;0;0;0m███[0m[38;2;15;0;0m█[0m[38;2;254;0;0m█[0m[38;2;252;0;0m█[0m[38;2;0;0;0m█[0m[38;2;0;2;0m█[0m[38;2;254;0;0m█[0m[38;2;254;0;2m█[0m[38;2;254;0;0m█[0m[38;2;254;5;1m█[0m[38;2;0;0;0m██[0m[38;2;174;14;16m█[0m[38;2;254;0;0m█[0m[38;2;255;5;0m█[0m[38;2;254;0;0m█[0m[38;2;32;0;0m█[0m[38;2;0;0;0m████████████████[0m[38;2;1;0;0m█[0m[38;2;122;85;69m█[0m[38;2;143;107;81m█[0m[38;2;176;145;125m█[0m[38;2;189;164;157m█[0m[38;2;187;164;150m█[0m[38;2;195;173;150m█[0m[38;2;188;172;156m█[0m[38;2;196;179;171m█[0m[38;2;201;183;179m█[0m[38;2;204;191;183m█[0m[38;2;197;188;183m█[0m[38;2;216;211;207m█[0m[38;2;239;235;232m█[0m[38;2;240;241;236m█[0m[38;2;237;239;234m█[0m[38;2;237;239;238m█[0m[38;2;240;239;244m█[0m[38;2;238;237;242m█[0m[38;2;241;241;241m█[0m[38;2;241;242;237m█[0m[38;2;239;240;235m█[0m[38;2;242;243;238m█[0m[38;2;240;241;236m█[0m[38;2;242;238;239m█[0m[38;2;241;237;234m█[0m[38;2;92;88;85m█[0m[38;2;165;159;163m█[0m[38;2;157;140;133m█[0m[38;2;190;173;155m█[0m[38;2;103;85;63m█[0m[38;2;84;62;38m█[0m[38;2;80;58;34m█[0m[38;2;109;83;56m█[0m[38;2;201;172;142m█[0m[38;2;207;175;137m█[0m[38;2;209;174;134m█[0m[38;2;224;185;142m█[0m[38;2;234;194;158m█[0m[38;2;235;200;162m█[0m[38;2;236;204;165m█[0m[38;2;231;202;158m█[0m[38;2;219;186;143m█[0m[38;2;210;176;141m█[0m[38;2;207;187;162m█[0m[38;2;30;29;25m█[0m[38;2;1;0;0m█[0m[38;2;0;0;0m███[0m");
$display("[38;2;0;0;0m████████████[0m[38;2;249;3;4m█[0m[38;2;254;0;0m█[0m[38;2;0;1;7m█[0m[38;2;0;0;0m███[0m[38;2;15;0;0m█[0m[38;2;254;0;0m█[0m[38;2;255;1;0m█[0m[38;2;0;0;0m█[0m[38;2;0;2;0m█[0m[38;2;254;0;0m█[0m[38;2;254;0;2m█[0m[38;2;129;0;0m█[0m[38;2;254;0;0m█[0m[38;2;29;0;0m█[0m[38;2;0;0;9m█[0m[38;2;251;2;0m█[0m[38;2;253;1;0m█[0m[38;2;255;1;1m█[0m[38;2;254;0;0m█[0m[38;2;32;0;0m█[0m[38;2;0;0;0m████████████████[0m[38;2;65;56;39m█[0m[38;2;138;111;84m█[0m[38;2;115;80;52m█[0m[38;2;162;131;113m█[0m[38;2;178;152;137m█[0m[38;2;180;152;140m█[0m[38;2;199;170;162m█[0m[38;2;210;193;186m█[0m[38;2;214;200;199m█[0m[38;2;222;213;214m█[0m[38;2;229;228;226m█[0m[38;2;231;230;228m█[0m[38;2;234;233;231m█[0m[38;2;235;235;235m█[0m[38;2;239;239;239m█[0m[38;2;240;240;240m██[0m[38;2;234;234;234m█[0m[38;2;241;241;241m███████[0m[38;2;235;235;235m█[0m[38;2;238;239;234m█[0m[38;2;145;145;135m█[0m[38;2;130;126;114m█[0m[38;2;85;79;63m█[0m[38;2;59;50;33m█[0m[38;2;192;177;156m█[0m[38;2;117;97;73m█[0m[38;2;198;177;146m█[0m[38;2;173;134;103m█[0m[38;2;191;146;113m█[0m[38;2;215;159;122m█[0m[38;2;229;177;137m█[0m[38;2;223;180;129m█[0m[38;2;221;180;128m█[0m[38;2;216;177;122m█[0m[38;2;207;173;128m█[0m[38;2;202;168;130m█[0m[38;2;199;168;137m█[0m[38;2;194;177;147m█[0m[38;2;89;85;73m█[0m[38;2;0;0;2m█[0m[38;2;0;0;0m███[0m");
$display("[38;2;0;0;0m████████████[0m[38;2;250;0;2m█[0m[38;2;254;0;0m█[0m[38;2;0;1;7m█[0m[38;2;0;0;0m███[0m[38;2;14;0;0m█[0m[38;2;254;0;0m█[0m[38;2;253;0;0m█[0m[38;2;0;0;0m█[0m[38;2;0;2;0m█[0m[38;2;254;0;0m█[0m[38;2;254;0;2m█[0m[38;2;0;0;2m█[0m[38;2;254;0;0m█[0m[38;2;255;4;4m█[0m[38;2;14;0;2m█[0m[38;2;253;1;0m█[0m[38;2;57;0;0m█[0m[38;2;255;2;0m█[0m[38;2;254;0;0m█[0m[38;2;32;0;0m█[0m[38;2;0;0;0m████████████████[0m[38;2;29;23;11m█[0m[38;2;129;92;83m█[0m[38;2;137;96;74m█[0m[38;2;155;123;108m█[0m[38;2;190;172;152m█[0m[38;2;189;176;159m█[0m[38;2;182;168;159m█[0m[38;2;213;200;192m█[0m[38;2;214;204;203m█[0m[38;2;209;198;204m█[0m[38;2;229;224;228m█[0m[38;2;218;213;217m█[0m[38;2;200;198;201m█[0m[38;2;224;224;224m█[0m[38;2;231;231;231m█[0m[38;2;241;241;241m███████████[0m[38;2;240;241;243m█[0m[38;2;238;238;238m█[0m[38;2;217;217;217m█[0m[38;2;175;175;173m█[0m[38;2;193;192;187m█[0m[38;2;177;173;162m█[0m[38;2;94;85;76m█[0m[38;2;102;81;62m█[0m[38;2;120;83;54m█[0m[38;2;187;146;118m█[0m[38;2;192;146;113m█[0m[38;2;203;157;121m█[0m[38;2;195;155;104m█[0m[38;2;208;161;119m█[0m[38;2;200;146;112m█[0m[38;2;191;144;102m█[0m[38;2;192;154;118m█[0m[38;2;191;162;132m█[0m[38;2;108;97;75m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m████████████[0m[38;2;254;1;0m█[0m[38;2;254;0;0m█[0m[38;2;166;15;6m█[0m[38;2;0;0;0m███[0m[38;2;237;18;12m█[0m[38;2;254;0;0m█[0m[38;2;241;2;5m█[0m[38;2;0;0;0m█[0m[38;2;0;2;0m█[0m[38;2;254;0;0m█[0m[38;2;254;0;2m█[0m[38;2;0;0;0m█[0m[38;2;218;16;12m█[0m[38;2;254;0;0m███[0m[38;2;0;1;2m█[0m[38;2;255;2;0m█[0m[38;2;254;0;0m█[0m[38;2;32;0;0m█[0m[38;2;0;0;0m████████████████[0m[38;2;1;0;0m█[0m[38;2;137;108;92m█[0m[38;2;112;78;53m█[0m[38;2;214;191;173m█[0m[38;2;192;170;157m█[0m[38;2;182;148;146m█[0m[38;2;179;169;160m█[0m[38;2;228;213;216m█[0m[38;2;222;212;210m█[0m[38;2;234;221;215m█[0m[38;2;223;215;212m█[0m[38;2;209;201;198m█[0m[38;2;183;180;175m█[0m[38;2;240;240;240m█[0m[38;2;242;242;242m██[0m[38;2;241;241;241m███████████[0m[38;2;242;242;242m█[0m[38;2;239;239;239m█[0m[38;2;236;236;238m█[0m[38;2;242;240;243m█[0m[38;2;227;222;219m█[0m[38;2;217;209;196m█[0m[38;2;184;166;152m█[0m[38;2;100;73;54m█[0m[38;2;91;59;34m█[0m[38;2;154;112;88m█[0m[38;2;158;104;78m█[0m[38;2;184;127;98m█[0m[38;2;172;119;85m█[0m[38;2;186;138;98m█[0m[38;2;195;147;111m█[0m[38;2;191;151;115m█[0m[38;2;180;154;117m█[0m[38;2;0;0;0m██████[0m");
$display("[38;2;0;0;0m████████████[0m[38;2;0;2;0m█[0m[38;2;249;0;9m█[0m[38;2;254;0;0m█████[0m[38;2;251;4;13m█[0m[38;2;1;0;0m█[0m[38;2;0;0;0m█[0m[38;2;0;2;0m█[0m[38;2;254;0;0m█[0m[38;2;254;0;2m█[0m[38;2;0;0;0m█[0m[38;2;0;1;4m█[0m[38;2;254;0;0m██[0m[38;2;102;0;0m█[0m[38;2;0;0;0m█[0m[38;2;255;2;0m█[0m[38;2;254;0;0m█[0m[38;2;32;0;0m█[0m[38;2;0;0;0m█[0m[38;2;1;0;0m█[0m[38;2;254;0;0m██[0m[38;2;0;0;0m███[0m[38;2;244;4;3m█[0m[38;2;254;0;0m█[0m[38;2;1;0;2m█[0m[38;2;0;0;0m█[0m[38;2;0;2;0m█[0m[38;2;254;0;0m█[0m[38;2;253;1;0m█[0m[38;2;0;0;0m██[0m[38;2;0;0;2m█[0m[38;2;102;96;74m█[0m[38;2;173;149;137m█[0m[38;2;222;205;197m█[0m[38;2;204;193;191m█[0m[38;2;208;197;193m█[0m[38;2;229;218;214m█[0m[38;2;228;220;217m██[0m[38;2;224;216;213m█[0m[38;2;225;217;214m█[0m[38;2;231;222;225m█[0m[38;2;247;238;241m█[0m[38;2;241;240;238m█[0m[38;2;242;241;239m█[0m[38;2;242;239;234m█[0m[38;2;239;240;235m██[0m[38;2;237;238;233m█[0m[38;2;239;239;237m█[0m[38;2;242;241;246m█[0m[38;2;241;241;241m████[0m[38;2;239;238;236m█[0m[38;2;232;228;225m█[0m[38;2;235;234;229m█[0m[38;2;239;241;238m█[0m[38;2;241;239;240m█[0m[38;2;238;237;235m█[0m[38;2;241;243;240m█[0m[38;2;237;239;234m█[0m[38;2;221;214;208m█[0m[38;2;118;97;94m█[0m[38;2;147;119;107m█[0m[38;2;84;66;46m█[0m[38;2;87;55;34m█[0m[38;2;149;99;76m█[0m[38;2;154;98;65m█[0m[38;2;167;121;95m█[0m[38;2;193;154;125m█[0m[38;2;183;150;115m█[0m[38;2;188;160;120m█[0m[38;2;63;56;38m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m██████████████[0m[38;2;0;1;0m█[0m[38;2;0;2;4m█[0m[38;2;3;0;4m█[0m[38;2;0;2;4m█[0m[38;2;0;1;0m█[0m[38;2;0;0;0m████████████████████████████████[0m[38;2;117;108;77m█[0m[38;2;234;232;237m█[0m[38;2;242;240;243m█[0m[38;2;241;241;239m██[0m[38;2;242;242;242m█[0m[38;2;238;237;242m█[0m[38;2;237;236;241m█[0m[38;2;228;227;225m█[0m[38;2;233;230;221m█[0m[38;2;235;225;216m█[0m[38;2;147;127;120m█[0m[38;2;79;51;37m█[0m[38;2;114;88;71m█[0m[38;2;137;111;96m█[0m[38;2;207;193;180m█[0m[38;2;207;208;194m█[0m[38;2;216;207;198m█[0m[38;2;235;227;224m█[0m[38;2;238;233;230m█[0m[38;2;241;241;241m███[0m[38;2;242;242;244m█[0m[38;2;220;205;202m█[0m[38;2;198;180;170m█[0m[38;2;194;182;170m█[0m[38;2;190;180;171m█[0m[38;2;200;186;185m█[0m[38;2;41;33;31m█[0m[38;2;44;36;34m█[0m[38;2;50;41;36m█[0m[38;2;86;71;66m█[0m[38;2;189;170;163m█[0m[38;2;88;80;69m█[0m[38;2;83;77;61m█[0m[38;2;118;102;86m█[0m[38;2;117;85;60m█[0m[38;2;146;105;73m█[0m[38;2;164;131;100m█[0m[38;2;172;143;113m█[0m[38;2;181;157;119m█[0m[38;2;74;62;48m█[0m[38;2;0;0;0m██████[0m");
$display("[38;2;0;0;0m██████████████████████████████████████████████████[0m[38;2;27;26;21m█[0m[38;2;242;229;223m█[0m[38;2;244;242;243m█[0m[38;2;244;239;243m█[0m[38;2;241;241;241m███[0m[38;2;242;241;246m█[0m[38;2;239;238;243m█[0m[38;2;242;237;241m█[0m[38;2;225;197;183m█[0m[38;2;180;146;119m█[0m[38;2;134;117;99m█[0m[38;2;76;80;79m█[0m[38;2;36;27;20m█[0m[38;2;152;120;79m█[0m[38;2;143;114;72m█[0m[38;2;174;146;135m█[0m[38;2;217;213;210m█[0m[38;2;228;227;225m█[0m[38;2;236;240;243m█[0m[38;2;241;241;241m██[0m[38;2;242;242;242m█[0m[38;2;233;232;228m█[0m[38;2;209;192;184m█[0m[38;2;194;170;158m█[0m[38;2;202;180;166m█[0m[38;2;45;28;10m█[0m[38;2;81;66;43m█[0m[38;2;92;86;72m█[0m[38;2;49;40;23m█[0m[38;2;98;78;53m█[0m[38;2;94;73;54m█[0m[38;2;60;44;31m█[0m[38;2;81;59;46m█[0m[38;2;71;54;46m█[0m[38;2;68;58;56m█[0m[38;2;96;78;76m█[0m[38;2;112;93;78m█[0m[38;2;77;55;42m█[0m[38;2;87;66;47m█[0m[38;2;142;126;101m█[0m[38;2;43;38;32m█[0m[38;2;0;0;0m██████[0m");
$display("[38;2;0;0;0m█████████████████████████████████████████████████[0m[38;2;74;75;69m█[0m[38;2;244;245;237m█[0m[38;2;241;241;239m█[0m[38;2;241;241;241m█████[0m[38;2;244;240;241m██[0m[38;2;245;241;240m█[0m[38;2;229;212;202m█[0m[38;2;200;179;152m█[0m[38;2;166;159;130m█[0m[38;2;39;36;29m█[0m[38;2;138;122;97m█[0m[38;2;191;168;118m█[0m[38;2;183;152;106m█[0m[38;2;131;109;98m█[0m[38;2;239;239;239m█[0m[38;2;241;241;241m████[0m[38;2;240;240;240m█[0m[38;2;240;238;239m█[0m[38;2;211;204;198m█[0m[38;2;212;200;188m█[0m[38;2;160;136;124m█[0m[38;2;118;93;73m█[0m[38;2;148;127;98m█[0m[38;2;73;71;58m█[0m[38;2;41;37;28m█[0m[38;2;86;66;41m█[0m[38;2;147;125;102m█[0m[38;2;70;47;29m█[0m[38;2;170;143;122m█[0m[38;2;158;140;126m█[0m[38;2;145;135;125m█[0m[38;2;71;66;62m█[0m[38;2;27;22;19m█[0m[38;2;64;58;60m█[0m[38;2;61;56;50m█[0m[38;2;82;80;59m█[0m[38;2;1;1;0m█[0m[38;2;0;0;0m██████[0m");
$display("[38;2;0;0;0m█████████████████████████████████████████████████[0m[38;2;233;231;216m█[0m[38;2;246;247;242m█[0m[38;2;240;240;240m█[0m[38;2;241;241;241m████[0m[38;2;242;240;241m█[0m[38;2;239;235;236m█[0m[38;2;242;238;239m█[0m[38;2;243;242;240m█[0m[38;2;238;238;240m█[0m[38;2;242;240;245m█[0m[38;2;252;243;238m█[0m[38;2;237;225;203m█[0m[38;2;222;219;204m█[0m[38;2;226;222;210m█[0m[38;2;244;230;227m█[0m[38;2;234;233;231m█[0m[38;2;240;242;241m█[0m[38;2;241;241;241m█████[0m[38;2;242;240;241m█[0m[38;2;247;241;243m█[0m[38;2;231;222;225m█[0m[38;2;200;195;189m█[0m[38;2;215;195;186m█[0m[38;2;76;54;33m█[0m[38;2;115;96;66m█[0m[38;2;122;106;80m█[0m[38;2;141;119;98m█[0m[38;2;170;153;143m█[0m[38;2;240;230;231m█[0m[38;2;217;213;214m█[0m[38;2;194;186;184m█[0m[38;2;138;128;126m█[0m[38;2;71;68;53m█[0m[38;2;117;113;104m█[0m[38;2;73;63;61m█[0m[38;2;63;44;48m█[0m[38;2;75;57;57m█[0m[38;2;64;51;45m█[0m[38;2;0;0;0m██████[0m");
$display("[38;2;0;0;0m████████████████████████████████████████████████[0m[38;2;19;18;16m█[0m[38;2;249;247;235m█[0m[38;2;245;238;245m█[0m[38;2;240;240;238m█[0m[38;2;241;241;241m█[0m[38;2;232;232;232m█[0m[38;2;233;235;234m█[0m[38;2;239;235;236m█[0m[38;2;228;222;224m█[0m[38;2;219;211;209m█[0m[38;2;218;210;208m█[0m[38;2;217;212;209m█[0m[38;2;232;232;232m█[0m[38;2;239;239;239m██[0m[38;2;241;241;239m██[0m[38;2;240;240;240m██[0m[38;2;241;241;241m█[0m[38;2;241;240;246m█[0m[38;2;241;240;245m██[0m[38;2;243;239;240m█[0m[38;2;242;238;239m██[0m[38;2;240;239;235m█[0m[38;2;230;226;223m█[0m[38;2;217;212;209m█[0m[38;2;233;233;235m█[0m[38;2;232;240;242m█[0m[38;2;234;239;242m█[0m[38;2;236;237;229m█[0m[38;2;237;238;232m█[0m[38;2;237;237;237m█[0m[38;2;226;227;221m█[0m[38;2;213;213;201m█[0m[38;2;201;201;191m█[0m[38;2;192;188;176m█[0m[38;2;190;181;166m█[0m[38;2;177;164;148m█[0m[38;2;172;158;149m█[0m[38;2;97;82;79m█[0m[38;2;71;55;55m█[0m[38;2;63;48;45m█[0m[38;2;59;44;39m█[0m[38;2;0;0;0m██████[0m");
$display("[38;2;0;0;0m█████████████████████████████████████████████████[0m[38;2;240;242;229m█[0m[38;2;241;241;241m█[0m[38;2;237;237;239m█[0m[38;2;233;233;233m█[0m[38;2;226;226;226m█[0m[38;2;225;229;232m█[0m[38;2;226;226;226m█[0m[38;2;206;205;201m█[0m[38;2;196;191;185m█[0m[38;2;191;186;182m█[0m[38;2;239;233;233m█[0m[38;2;239;235;236m█[0m[38;2;243;239;240m█[0m[38;2;241;237;238m██[0m[38;2;241;239;242m█[0m[38;2;240;244;245m█[0m[38;2;243;243;245m█[0m[38;2;232;230;233m█[0m[38;2;239;234;230m█[0m[38;2;245;229;229m█[0m[38;2;233;211;213m█[0m[38;2;221;191;191m█[0m[38;2;226;197;193m█[0m[38;2;223;194;186m█[0m[38;2;202;170;157m█[0m[38;2;209;171;162m█[0m[38;2;207;169;160m█[0m[38;2;181;157;155m█[0m[38;2;200;196;197m█[0m[38;2;214;205;210m█[0m[38;2;212;201;207m█[0m[38;2;205;196;191m█[0m[38;2;195;196;191m█[0m[38;2;202;199;194m█[0m[38;2;200;186;183m█[0m[38;2;189;175;164m█[0m[38;2;167;149;135m█[0m[38;2;177;154;136m█[0m[38;2;174;156;134m█[0m[38;2;178;159;142m█[0m[38;2;165;146;132m█[0m[38;2;63;46;36m█[0m[38;2;54;41;33m█[0m[38;2;63;52;48m█[0m[38;2;172;158;158m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m████████████████████████████████████████████████[0m[38;2;170;170;168m█[0m[38;2;238;238;236m█[0m[38;2;240;241;236m█[0m[38;2;226;226;224m█[0m[38;2;223;223;223m█[0m[38;2;224;224;224m█[0m[38;2;229;225;222m█[0m[38;2;203;196;190m█[0m[38;2;187;176;170m█[0m[38;2;188;175;169m█[0m[38;2;228;227;222m█[0m[38;2;221;221;219m█[0m[38;2;203;192;196m█[0m[38;2;200;189;193m█[0m[38;2;196;186;187m█[0m[38;2;233;224;219m█[0m[38;2;218;209;204m█[0m[38;2;209;206;199m█[0m[38;2;212;207;201m█[0m[38;2;228;217;213m█[0m[38;2;227;196;202m█[0m[38;2;204;159;156m█[0m[38;2;196;133;128m█[0m[38;2;183;114;98m█[0m[38;2;181;113;92m█[0m[38;2;177;111;85m█[0m[38;2;157;91;77m█[0m[38;2;141;83;69m█[0m[38;2;190;144;128m█[0m[38;2;187;163;151m█[0m[38;2;187;169;165m█[0m[38;2;185;166;160m█[0m[38;2;181;166;159m█[0m[38;2;184;169;164m█[0m[38;2;189;174;169m█[0m[38;2;191;178;169m█[0m[38;2;191;182;165m█[0m[38;2;195;178;168m█[0m[38;2;193;175;161m█[0m[38;2;175;152;134m█[0m[38;2;163;146;118m█[0m[38;2;166;148;124m█[0m[38;2;177;159;137m█[0m[38;2;155;134;115m█[0m[38;2;98;81;65m█[0m[38;2;97;81;66m█[0m[38;2;171;157;144m█[0m[38;2;79;76;69m█[0m[38;2;0;1;0m█[0m[38;2;0;0;0m███[0m");
$display("[38;2;0;0;0m█████████████████████████████████████████████[0m[38;2;61;60;58m█[0m[38;2;232;228;225m█[0m[38;2;240;240;242m█[0m[38;2;243;243;243m█[0m[38;2;242;242;242m█[0m[38;2;240;240;240m█[0m[38;2;227;228;230m█[0m[38;2;223;222;220m█[0m[38;2;217;210;204m█[0m[38;2;204;199;195m█[0m[38;2;196;187;180m█[0m[38;2;202;192;182m█[0m[38;2;208;203;199m█[0m[38;2;213;208;204m█[0m[38;2;192;189;184m█[0m[38;2;165;164;159m█[0m[38;2;176;168;165m█[0m[38;2;173;163;161m█[0m[38;2;164;153;147m█[0m[38;2;166;156;146m█[0m[38;2;173;163;151m█[0m[38;2;174;161;152m█[0m[38;2;173;156;148m█[0m[38;2;157;151;127m█[0m[38;2;161;149;123m█[0m[38;2;172;136;114m█[0m[38;2;170;118;96m█[0m[38;2;154;97;78m█[0m[38;2;154;96;76m█[0m[38;2;157;119;100m█[0m[38;2;149;126;110m█[0m[38;2;154;137;121m█[0m[38;2;156;135;118m█[0m[38;2;168;147;130m█[0m[38;2;169;147;134m█[0m[38;2;166;144;133m█[0m[38;2;156;134;123m█[0m[38;2;159;136;122m█[0m[38;2;153;130;114m█[0m[38;2;156;134;111m█[0m[38;2;162;139;123m█[0m[38;2;176;153;137m█[0m[38;2;179;156;140m█[0m[38;2;176;154;140m█[0m[38;2;178;151;140m█[0m[38;2;178;150;136m█[0m[38;2;182;154;140m█[0m[38;2;174;151;135m█[0m[38;2;170;153;135m█[0m[38;2;191;179;165m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m██████████████████████████████████████████[0m[38;2;22;22;20m█[0m[38;2;122;123;115m█[0m[38;2;235;235;233m█[0m[38;2;244;244;246m█[0m[38;2;242;242;242m█[0m[38;2;241;241;241m███[0m[38;2;244;244;244m█[0m[38;2;232;226;230m█[0m[38;2;224;220;219m█[0m[38;2;213;210;203m█[0m[38;2;209;202;196m█[0m[38;2;203;193;184m█[0m[38;2;199;185;174m█[0m[38;2;189;181;170m█[0m[38;2;185;177;166m█[0m[38;2;177;168;159m█[0m[38;2;164;155;148m█[0m[38;2;155;142;133m█[0m[38;2;138;124;111m█[0m[38;2;117;99;85m█[0m[38;2;116;94;81m█[0m[38;2;114;95;81m█[0m[38;2;126;104;91m█[0m[38;2;136;109;98m█[0m[38;2;133;109;105m█[0m[38;2;138;109;101m█[0m[38;2;138;105;96m█[0m[38;2;132;92;84m█[0m[38;2;127;82;76m█[0m[38;2;121;81;73m█[0m[38;2;122;88;87m█[0m[38;2;130;102;99m██[0m[38;2;126;97;91m█[0m[38;2;122;94;83m█[0m[38;2;120;92;81m█[0m[38;2;118;90;79m█[0m[38;2;117;89;78m█[0m[38;2;122;96;79m█[0m[38;2;154;129;107m█[0m[38;2;158;134;108m█[0m[38;2;162;136;121m█[0m[38;2;161;135;118m█[0m[38;2;164;138;121m█[0m[38;2;164;140;116m█[0m[38;2;170;146;122m█[0m[38;2;178;153;131m█[0m[38;2;180;152;140m█[0m[38;2;176;154;131m█[0m[38;2;170;152;128m█[0m[38;2;157;145;131m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m█████████████████████████████████████████[0m[38;2;167;166;171m█[0m[38;2;249;248;254m█[0m[38;2;241;240;245m█[0m[38;2;241;241;243m█[0m[38;2;241;241;241m██████[0m[38;2;236;230;234m█[0m[38;2;231;227;226m█[0m[38;2;227;224;217m█[0m[38;2;203;196;190m█[0m[38;2;198;188;179m█[0m[38;2;197;183;172m█[0m[38;2;188;180;169m█[0m[38;2;181;173;162m█[0m[38;2;175;166;157m█[0m[38;2;168;159;152m█[0m[38;2;164;151;142m█[0m[38;2;156;142;129m█[0m[38;2;148;132;117m█[0m[38;2;141;119;106m█[0m[38;2;145;126;112m█[0m[38;2;148;126;113m█[0m[38;2;144;117;106m█[0m[38;2;137;115;101m█[0m[38;2;133;105;91m█[0m[38;2;128;97;79m█[0m[38;2;120;94;81m█[0m[38;2;136;99;90m█[0m[38;2;140;99;93m█[0m[38;2;130;97;88m█[0m[38;2;132;105;94m█[0m[38;2;131;104;97m█[0m[38;2;136;107;101m█[0m[38;2;138;110;99m█[0m[38;2;139;111;97m█[0m[38;2;137;110;91m█[0m[38;2;139;112;93m█[0m[38;2;140;114;97m█[0m[38;2;146;121;99m█[0m[38;2;155;131;105m█[0m[38;2;158;134;108m█[0m[38;2;162;138;112m█[0m[38;2;166;142;116m█[0m[38;2;170;146;122m█[0m[38;2;171;147;123m█[0m[38;2;169;148;121m█[0m[38;2;170;150;125m█[0m[38;2;169;152;132m█[0m[38;2;172;159;143m█[0m[38;2;89;82;72m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m███████████████████████████████████████[0m[38;2;31;31;33m█[0m[38;2;229;229;229m█[0m[38;2;241;241;241m█[0m[38;2;243;243;243m█[0m[38;2;241;241;241m████████[0m[38;2;231;231;229m█[0m[38;2;225;224;219m█[0m[38;2;205;201;192m█[0m[38;2;198;190;179m█[0m[38;2;195;187;176m█[0m[38;2;191;183;172m█[0m[38;2;188;180;169m█[0m[38;2;180;172;161m█[0m[38;2;176;166;156m█[0m[38;2;169;155;146m█[0m[38;2;171;158;142m█[0m[38;2;164;151;134m█[0m[38;2;169;153;138m█[0m[38;2;163;146;136m█[0m[38;2;161;147;134m█[0m[38;2;160;147;131m█[0m[38;2;151;138;122m█[0m[38;2;152;134;124m█[0m[38;2;154;131;125m█[0m[38;2;154;125;119m█[0m[38;2;152;126;111m█[0m[38;2;149;123;108m█[0m[38;2;152;126;111m█[0m[38;2;155;127;113m█[0m[38;2;149;126;110m█[0m[38;2;154;131;117m█[0m[38;2;152;126;113m█[0m[38;2;149;123;106m█[0m[38;2;154;129;107m█[0m[38;2;150;125;103m█[0m[38;2;152;127;105m█[0m[38;2;155;131;107m█[0m[38;2;158;134;110m█[0m[38;2;162;138;114m██[0m[38;2;164;140;116m█[0m[38;2;168;144;120m█[0m[38;2;170;146;122m█[0m[38;2;171;147;123m█[0m[38;2;174;150;126m█[0m[38;2;172;152;127m█[0m[38;2;173;156;136m█[0m[38;2;191;178;161m█[0m[38;2;11;10;8m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m██████████████████████████████████████[0m[38;2;119;118;123m█[0m[38;2;230;229;234m█[0m[38;2;241;241;239m█[0m[38;2;242;242;242m██[0m[38;2;241;241;241m████████[0m[38;2;240;238;241m█[0m[38;2;238;232;232m█[0m[38;2;223;214;209m█[0m[38;2;209;200;191m█[0m[38;2;194;185;176m█[0m[38;2;191;182;173m█[0m[38;2;183;174;169m█[0m[38;2;178;169;160m█[0m[38;2;178;170;157m█[0m[38;2;174;164;152m█[0m[38;2;175;159;144m█[0m[38;2;173;157;141m█[0m[38;2;169;156;140m█[0m[38;2;162;149;133m█[0m[38;2;156;147;130m█[0m[38;2;156;149;131m█[0m[38;2;155;148;130m█[0m[38;2;151;140;120m█[0m[38;2;151;136;117m█[0m[38;2;153;136;118m█[0m[38;2;152;129;113m█[0m[38;2;155;127;113m█[0m[38;2;156;127;113m█[0m[38;2;156;126;118m█[0m[38;2;156;126;116m█[0m[38;2;154;127;116m█[0m[38;2;150;131;114m█[0m[38;2;149;131;109m█[0m[38;2;152;131;110m█[0m[38;2;152;134;110m█[0m[38;2;153;136;106m█[0m[38;2;161;135;98m█[0m[38;2;166;140;105m█[0m[38;2;167;140;110m█[0m[38;2;167;138;124m█[0m[38;2;173;144;128m██[0m[38;2;171;147;123m█[0m[38;2;173;149;125m█[0m[38;2;178;154;130m█[0m[38;2;171;151;126m█[0m[38;2;174;157;137m█[0m[38;2;195;182;165m█[0m[38;2;0;0;0m██████[0m");
$display("[38;2;0;0;0m████████████████████████████████████[0m[38;2;3;3;3m█[0m[38;2;196;195;200m█[0m[38;2;238;237;242m█[0m[38;2;241;240;245m█[0m[38;2;241;241;239m█[0m[38;2;241;241;241m██████████[0m[38;2;241;239;242m█[0m[38;2;236;230;230m█[0m[38;2;222;213;208m█[0m[38;2;200;191;182m█[0m[38;2;194;185;176m█[0m[38;2;189;180;171m█[0m[38;2;182;173;168m█[0m[38;2;179;170;161m█[0m[38;2;178;170;157m█[0m[38;2;179;169;157m█[0m[38;2;180;164;149m█[0m[38;2;175;159;143m█[0m[38;2;168;155;139m█[0m[38;2;164;151;135m█[0m[38;2;163;148;127m█[0m[38;2;160;145;122m█[0m[38;2;163;148;125m█[0m[38;2;157;146;126m█[0m[38;2;156;141;122m█[0m[38;2;158;139;122m█[0m[38;2;149;134;115m█[0m[38;2;146;127;110m█[0m[38;2;154;133;116m█[0m[38;2;154;134;110m█[0m[38;2;151;130;109m█[0m[38;2;149;131;111m█[0m[38;2;152;134;110m█[0m[38;2;151;134;106m█[0m[38;2;156;134;110m█[0m[38;2;165;138;117m█[0m[38;2;163;137;110m█[0m[38;2;160;141;108m█[0m[38;2;164;145;115m█[0m[38;2;164;144;119m█[0m[38;2;167;147;120m█[0m[38;2;168;148;123m██[0m[38;2;171;147;123m██[0m[38;2;174;150;126m█[0m[38;2;174;153;136m█[0m[38;2;189;171;157m█[0m[38;2;213;201;189m█[0m[38;2;56;52;49m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m███████████████████████████████████[0m[38;2;76;74;77m█[0m[38;2;200;195;202m█[0m[38;2;242;242;242m█[0m[38;2;241;241;241m█████████████[0m[38;2;240;238;241m█[0m[38;2;241;235;235m█[0m[38;2;231;221;219m█[0m[38;2;210;210;202m█[0m[38;2;190;186;175m█[0m[38;2;188;180;167m█[0m[38;2;183;174;169m█[0m[38;2;180;171;162m█[0m[38;2;180;172;159m█[0m[38;2;178;169;152m█[0m[38;2;183;167;152m█[0m[38;2;180;164;149m█[0m[38;2;173;161;139m█[0m[38;2;170;157;138m█[0m[38;2;164;156;135m█[0m[38;2;158;147;127m█[0m[38;2;163;148;129m█[0m[38;2;161;146;127m█[0m[38;2;156;141;122m█[0m[38;2;152;137;118m█[0m[38;2;154;136;114m█[0m[38;2;151;133;111m██[0m[38;2;153;135;113m█[0m[38;2;152;134;112m█[0m[38;2;151;133;109m█[0m[38;2;156;139;113m██[0m[38;2;160;143;117m█[0m[38;2;163;146;120m█[0m[38;2;167;143;119m█[0m[38;2;167;145;121m█[0m[38;2;166;146;121m█[0m[38;2;165;145;120m█[0m[38;2;168;148;123m█[0m[38;2;168;148;121m█[0m[38;2;168;149;117m█[0m[38;2;173;149;123m█[0m[38;2;173;148;126m█[0m[38;2;178;152;135m█[0m[38;2;179;160;143m█[0m[38;2;190;173;166m█[0m[38;2;201;187;187m█[0m[38;2;154;146;143m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m██████████████████████████████████[0m[38;2;133;131;142m█[0m[38;2;167;166;172m█[0m[38;2;232;232;234m█[0m[38;2;242;242;242m██[0m[38;2;241;241;241m███████████[0m[38;2;238;238;238m█[0m[38;2;238;239;241m█[0m[38;2;239;238;236m█[0m[38;2;229;224;218m█[0m[38;2;208;201;195m█[0m[38;2;197;187;178m█[0m[38;2;193;179;168m█[0m[38;2;178;169;164m█[0m[38;2;177;168;159m█[0m[38;2;173;165;152m█[0m[38;2;174;165;148m█[0m[38;2;177;161;146m█[0m[38;2;178;160;146m█[0m[38;2;169;160;143m█[0m[38;2;166;157;140m█[0m[38;2;163;156;137m█[0m[38;2;162;151;131m█[0m[38;2;160;145;126m█[0m[38;2;159;142;124m█[0m[38;2;159;140;123m█[0m[38;2;160;137;121m█[0m[38;2;157;140;112m█[0m[38;2;153;136;110m█[0m[38;2;153;135;115m██[0m[38;2;152;135;109m█[0m[38;2;156;139;113m█[0m[38;2;157;140;114m█[0m[38;2;160;143;117m█[0m[38;2;162;144;122m█[0m[38;2;166;149;123m█[0m[38;2;166;146;119m█[0m[38;2;166;146;122m█[0m[38;2;169;144;122m█[0m[38;2;172;143;127m█[0m[38;2;171;145;122m█[0m[38;2;170;145;125m█[0m[38;2;170;144;127m█[0m[38;2;171;147;123m█[0m[38;2;178;154;130m█[0m[38;2;185;161;135m█[0m[38;2;188;163;141m█[0m[38;2;193;174;157m█[0m[38;2;204;186;172m█[0m[38;2;145;133;117m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m█████████████████████████████████[0m[38;2;15;15;17m█[0m[38;2;199;197;210m█[0m[38;2;238;237;243m█[0m[38;2;243;243;245m█[0m[38;2;242;242;242m██[0m[38;2;241;241;241m████████████[0m[38;2;236;237;239m█[0m[38;2;226;225;223m█[0m[38;2;214;209;203m█[0m[38;2;220;213;207m█[0m[38;2;207;197;188m█[0m[38;2;198;184;173m█[0m[38;2;183;174;169m█[0m[38;2;178;169;160m█[0m[38;2;174;166;153m█[0m[38;2;168;159;142m█[0m[38;2;172;156;141m█[0m[38;2;170;154;139m█[0m[38;2;165;156;139m█[0m[38;2;163;154;137m█[0m[38;2;161;154;135m█[0m[38;2;162;151;131m█[0m[38;2;165;150;131m█[0m[38;2;158;147;127m█[0m[38;2;161;146;127m█[0m[38;2;162;143;126m█[0m[38;2;160;143;117m█[0m[38;2;156;140;107m█[0m[38;2;160;144;111m█[0m[38;2;158;142;109m█[0m[38;2;157;140;112m█[0m[38;2;157;140;114m█[0m[38;2;158;141;115m█[0m[38;2;159;142;116m█[0m[38;2;160;142;120m█[0m[38;2;165;147;123m█[0m[38;2;162;145;115m█[0m[38;2;158;143;112m█[0m[38;2;159;144;113m█[0m[38;2;162;143;113m█[0m[38;2;165;142;111m█[0m[38;2;167;143;115m█[0m[38;2;170;146;122m█[0m[38;2;174;150;126m█[0m[38;2;180;156;132m█[0m[38;2;185;161;135m█[0m[38;2;190;165;145m█[0m[38;2;193;172;155m█[0m[38;2;199;181;167m█[0m[38;2;165;153;141m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m████████████████████████████████[0m[38;2;0;0;2m█[0m[38;2;176;175;181m█[0m[38;2;221;219;230m█[0m[38;2;246;245;251m█[0m[38;2;239;239;241m█[0m[38;2;242;242;242m██[0m[38;2;241;241;241m███████████[0m[38;2;238;238;238m█[0m[38;2;234;233;231m█[0m[38;2;235;230;227m█[0m[38;2;225;216;211m█[0m[38;2;211;210;206m█[0m[38;2;207;203;194m█[0m[38;2;202;194;183m█[0m[38;2;189;180;175m█[0m[38;2;185;176;167m█[0m[38;2;180;173;157m█[0m[38;2;172;164;143m█[0m[38;2;168;160;139m█[0m[38;2;167;159;138m█[0m[38;2;162;154;133m█[0m[38;2;162;149;130m█[0m[38;2;164;147;127m█[0m[38;2;161;149;127m█[0m[38;2;159;151;128m█[0m[38;2;163;150;131m█[0m[38;2;165;150;131m█[0m[38;2;167;148;131m█[0m[38;2;157;140;114m█[0m[38;2;160;143;117m███[0m[38;2;157;140;114m██[0m[38;2;158;141;115m██[0m[38;2;156;138;116m█[0m[38;2;161;143;119m█[0m[38;2;161;144;114m█[0m[38;2;162;142;115m██[0m[38;2;162;142;117m█[0m[38;2;173;144;114m█[0m[38;2;171;146;116m█[0m[38;2;172;150;126m█[0m[38;2;175;155;128m█[0m[38;2;181;156;134m█[0m[38;2;188;161;144m█[0m[38;2;186;168;146m█[0m[38;2;187;172;153m█[0m[38;2;196;184;168m█[0m[38;2;201;193;172m█[0m[38;2;185;177;154m█[0m[38;2;1;0;0m█[0m[38;2;0;0;0m███[0m");
$display("[38;2;0;0;0m███████████████████████████████[0m[38;2;99;98;103m█[0m[38;2;161;160;168m█[0m[38;2;211;210;218m█[0m[38;2;240;239;245m█[0m[38;2;242;241;246m█[0m[38;2;241;241;241m█████████████[0m[38;2;233;233;233m█[0m[38;2;230;230;230m█[0m[38;2;228;228;230m█[0m[38;2;223;219;220m█[0m[38;2;221;213;211m█[0m[38;2;219;215;212m█[0m[38;2;208;201;195m█[0m[38;2;206;196;187m█[0m[38;2;193;184;179m█[0m[38;2;188;179;170m█[0m[38;2;183;176;160m█[0m[38;2;178;172;150m█[0m[38;2;174;166;145m█[0m[38;2;171;163;142m█[0m[38;2;176;163;146m█[0m[38;2;177;161;145m█[0m[38;2;179;156;140m█[0m[38;2;176;155;138m█[0m[38;2;170;153;135m█[0m[38;2;172;151;134m█[0m[38;2;167;146;129m█[0m[38;2;167;144;128m█[0m[38;2;164;148;125m█[0m[38;2;154;136;112m█[0m[38;2;166;142;116m█[0m[38;2;160;142;118m█[0m[38;2;158;141;115m█[0m[38;2;158;141;113m█[0m[38;2;160;143;115m█[0m[38;2;161;144;118m█[0m[38;2;159;141;117m█[0m[38;2;163;145;123m█[0m[38;2;164;147;119m█[0m[38;2;171;146;116m█[0m[38;2;171;144;115m█[0m[38;2;171;146;115m█[0m[38;2;170;150;113m█[0m[38;2;169;153;120m█[0m[38;2;170;156;127m█[0m[38;2;177;156;129m█[0m[38;2;179;155;131m█[0m[38;2;188;161;142m█[0m[38;2;185;163;142m█[0m[38;2;187;166;149m█[0m[38;2;196;177;163m█[0m[38;2;203;187;174m█[0m[38;2;211;194;178m█[0m[38;2;0;0;2m█[0m[38;2;0;0;0m███[0m");
$display("[38;2;0;0;0m██████████████████████████████[0m[38;2;102;101;106m█[0m[38;2;174;173;179m█[0m[38;2;213;212;218m█[0m[38;2;242;241;247m█[0m[38;2;241;241;241m██████████████[0m[38;2;239;239;239m█[0m[38;2;234;234;234m█[0m[38;2;225;225;225m█[0m[38;2;215;216;218m█[0m[38;2;220;219;217m█[0m[38;2;221;214;208m█[0m[38;2;211;211;209m█[0m[38;2;207;204;199m█[0m[38;2;204;197;187m█[0m[38;2;196;187;182m█[0m[38;2;194;185;176m█[0m[38;2;189;181;168m█[0m[38;2;186;179;163m█[0m[38;2;178;171;155m█[0m[38;2;174;167;151m█[0m[38;2;174;165;148m█[0m[38;2;172;163;146m█[0m[38;2;171;158;139m█[0m[38;2;173;158;139m██[0m[38;2;169;154;135m██[0m[38;2;166;153;134m█[0m[38;2;166;149;129m█[0m[38;2;167;147;123m█[0m[38;2;170;146;120m█[0m[38;2;166;148;124m█[0m[38;2;163;146;120m█[0m[38;2;159;142;114m█[0m[38;2;160;143;113m█[0m[38;2;158;141;115m█[0m[38;2;160;139;118m█[0m[38;2;166;145;124m█[0m[38;2;166;146;119m█[0m[38;2;167;144;113m█[0m[38;2;170;147;116m█[0m[38;2;175;152;121m█[0m[38;2;173;150;119m█[0m[38;2;175;151;127m█[0m[38;2;176;149;130m█[0m[38;2;182;158;134m█[0m[38;2;181;157;133m██[0m[38;2;184;159;137m█[0m[38;2;186;165;146m█[0m[38;2;189;173;157m█[0m[38;2;187;174;157m█[0m[38;2;0;1;0m█[0m[38;2;1;0;0m█[0m[38;2;0;0;0m███[0m");
$display("[38;2;0;0;0m████████████████████████████[0m[38;2;24;24;22m█[0m[38;2;168;169;161m█[0m[38;2;175;174;180m█[0m[38;2;189;187;198m█[0m[38;2;235;234;239m█[0m[38;2;243;243;243m█[0m[38;2;241;241;241m██████████████[0m[38;2;242;242;242m█[0m[38;2;236;236;236m█[0m[38;2;232;232;234m█[0m[38;2;229;228;233m█[0m[38;2;219;219;219m█[0m[38;2;219;220;215m█[0m[38;2;215;214;212m█[0m[38;2;211;206;202m█[0m[38;2;208;199;192m█[0m[38;2;203;194;185m█[0m[38;2;198;189;180m█[0m[38;2;189;180;171m█[0m[38;2;186;175;169m█[0m[38;2;184;174;164m█[0m[38;2;179;170;155m█[0m[38;2;181;168;152m█[0m[38;2;180;167;151m█[0m[38;2;176;163;147m██[0m[38;2;174;161;145m█[0m[38;2;170;165;136m█[0m[38;2;168;158;133m█[0m[38;2;173;157;141m█[0m[38;2;170;158;142m█[0m[38;2;167;152;133m█[0m[38;2;165;147;125m█[0m[38;2;171;153;129m█[0m[38;2;167;149;125m█[0m[38;2;163;149;123m█[0m[38;2;164;153;125m█[0m[38;2;169;149;124m█[0m[38;2;168;144;120m██[0m[38;2;169;145;121m█[0m[38;2;167;143;119m█[0m[38;2;170;146;118m█[0m[38;2;172;149;117m█[0m[38;2;174;149;119m█[0m[38;2;176;150;125m█[0m[38;2;177;150;131m█[0m[38;2;175;158;132m█[0m[38;2;180;156;132m█[0m[38;2;181;155;132m█[0m[38;2;183;159;133m█[0m[38;2;184;164;140m█[0m[38;2;184;167;149m█[0m[38;2;191;175;160m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m███████████████████████████[0m[38;2;3;3;3m█[0m[38;2;156;146;154m█[0m[38;2;179;178;184m█[0m[38;2;200;199;205m█[0m[38;2;228;227;235m█[0m[38;2;241;240;246m█[0m[38;2;242;242;242m█[0m[38;2;241;241;241m██████████████[0m[38;2;239;239;239m█[0m[38;2;234;234;234m█[0m[38;2;228;228;226m█[0m[38;2;217;218;212m█[0m[38;2;216;219;210m█[0m[38;2;213;215;202m█[0m[38;2;209;208;206m█[0m[38;2;208;203;199m█[0m[38;2;203;194;187m█[0m[38;2;199;190;181m█[0m[38;2;198;189;180m█[0m[38;2;190;181;172m█[0m[38;2;189;178;172m█[0m[38;2;184;174;164m█[0m[38;2;184;172;158m█[0m[38;2;181;169;153m█[0m[38;2;179;167;151m█[0m[38;2;178;165;149m█[0m[38;2;175;162;146m█[0m[38;2;177;164;148m█[0m[38;2;168;161;145m█[0m[38;2;171;160;138m█[0m[38;2;174;159;128m█[0m[38;2;173;161;145m█[0m[38;2;172;159;140m█[0m[38;2;172;156;131m█[0m[38;2;166;152;126m█[0m[38;2;168;150;126m█[0m[38;2;165;148;120m█[0m[38;2;166;149;123m█[0m[38;2;162;146;120m█[0m[38;2;166;149;121m█[0m[38;2;169;147;123m█[0m[38;2;169;147;124m█[0m[38;2;167;145;122m█[0m[38;2;172;151;120m█[0m[38;2;175;150;120m█[0m[38;2;170;154;121m█[0m[38;2;174;154;127m█[0m[38;2;174;156;134m█[0m[38;2;178;158;133m█[0m[38;2;181;157;133m█[0m[38;2;182;156;133m█[0m[38;2;178;156;132m█[0m[38;2;181;160;139m█[0m[38;2;183;166;148m█[0m[38;2;136;124;110m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m██████████████████████████[0m[38;2;14;15;10m█[0m[38;2;180;185;163m█[0m[38;2;181;186;182m█[0m[38;2;184;183;189m█[0m[38;2;196;195;201m█[0m[38;2;225;225;227m█[0m[38;2;241;241;241m██████[0m[38;2;240;240;240m█[0m[38;2;242;242;242m██[0m[38;2;240;240;240m█[0m[38;2;241;241;241m█[0m[38;2;237;237;237m█[0m[38;2;241;241;241m█[0m[38;2;242;242;242m█[0m[38;2;241;241;243m█[0m[38;2;244;243;249m█[0m[38;2;235;235;243m█[0m[38;2;232;230;235m█[0m[38;2;232;226;228m█[0m[38;2;219;218;216m█[0m[38;2;216;213;208m█[0m[38;2;207;204;195m█[0m[38;2;207;202;196m█[0m[38;2;209;204;198m█[0m[38;2;206;201;195m█[0m[38;2;194;195;181m█[0m[38;2;189;185;173m█[0m[38;2;193;184;175m█[0m[38;2;184;175;168m█[0m[38;2;186;178;167m█[0m[38;2;182;173;158m█[0m[38;2;177;165;149m██[0m[38;2;181;168;152m█[0m[38;2;181;168;149m█[0m[38;2;177;165;143m█[0m[38;2;167;160;142m█[0m[38;2;170;159;139m█[0m[38;2;174;159;136m█[0m[38;2;172;159;143m█[0m[38;2;173;160;141m█[0m[38;2;168;156;132m█[0m[38;2;168;151;125m█[0m[38;2;168;150;126m█[0m[38;2;169;151;127m█[0m[38;2;169;152;126m██[0m[38;2;171;151;126m█[0m[38;2;171;149;125m█[0m[38;2;167;146;117m█[0m[38;2;167;146;115m██[0m[38;2;170;149;118m█[0m[38;2;167;148;116m█[0m[38;2;168;144;120m█[0m[38;2;174;145;127m█[0m[38;2;179;155;131m█[0m[38;2;181;157;133m█[0m[38;2;178;156;132m█[0m[38;2;183;156;135m█[0m[38;2;180;158;135m█[0m[38;2;180;162;142m█[0m[38;2;128;114;101m█[0m[38;2;0;0;0m█████[0m");
$display("[38;2;0;0;0m█████████████████████████[0m[38;2;1;1;1m█[0m[38;2;115;106;89m█[0m[38;2;170;170;160m█[0m[38;2;171;174;179m█[0m[38;2;178;177;183m█[0m[38;2;213;212;218m█[0m[38;2;241;241;243m█[0m[38;2;241;241;241m█████[0m[38;2;236;236;236m█[0m[38;2;234;234;234m█[0m[38;2;238;238;238m█[0m[38;2;236;236;236m█[0m[38;2;229;229;229m█[0m[38;2;226;226;226m█[0m[38;2;230;230;230m█[0m[38;2;234;234;234m█[0m[38;2;238;238;238m█[0m[38;2;237;237;237m█[0m[38;2;238;237;243m█[0m[38;2;230;231;233m█[0m[38;2;227;225;226m█[0m[38;2;223;217;221m█[0m[38;2;213;207;207m█[0m[38;2;209;204;200m█[0m[38;2;212;208;199m█[0m[38;2;207;202;196m█[0m[38;2;198;193;187m██[0m[38;2;202;193;186m█[0m[38;2;200;191;182m█[0m[38;2;199;191;180m█[0m[38;2;189;179;170m█[0m[38;2;186;177;160m█[0m[38;2;184;176;157m█[0m[38;2;184;172;148m█[0m[38;2;180;168;144m█[0m[38;2;175;163;139m█[0m[38;2;175;160;137m█[0m[38;2;173;158;135m█[0m[38;2;171;163;144m█[0m[38;2;169;162;136m█[0m[38;2;168;161;132m█[0m[38;2;164;156;135m█[0m[38;2;172;160;136m█[0m[38;2;175;159;133m█[0m[38;2;176;154;130m█[0m[38;2;174;150;126m█[0m[38;2;176;154;130m█[0m[38;2;172;155;129m█[0m[38;2;169;152;126m█[0m[38;2;167;149;127m█[0m[38;2;167;149;125m█[0m[38;2;171;150;121m█[0m[38;2;174;151;120m█[0m[38;2;170;147;116m█[0m[38;2;172;149;118m█[0m[38;2;175;151;127m█[0m[38;2;176;152;128m██[0m[38;2;175;149;122m█[0m[38;2;174;148;121m██[0m[38;2;176;151;129m█[0m[38;2;173;152;135m█[0m[38;2;176;159;143m█[0m[38;2;0;0;0m██████[0m");
$display("[38;2;0;0;0m█████████████████████████[0m[38;2;1;1;1m█[0m[38;2;125;123;110m█[0m[38;2;169;164;161m█[0m[38;2;149;136;153m█[0m[38;2;181;182;186m█[0m[38;2;226;225;231m█[0m[38;2;242;242;242m██[0m[38;2;241;241;241m█[0m[38;2;242;242;242m██[0m[38;2;238;238;238m█[0m[38;2;233;233;233m█[0m[38;2;231;231;231m██[0m[38;2;228;228;228m█[0m[38;2;224;224;224m█[0m[38;2;219;219;219m█[0m[38;2;215;215;215m█[0m[38;2;223;223;223m█[0m[38;2;224;224;224m█[0m[38;2;228;228;230m█[0m[38;2;226;225;233m█[0m[38;2;220;222;217m█[0m[38;2;213;214;206m█[0m[38;2;212;209;202m█[0m[38;2;200;196;195m█[0m[38;2;206;203;198m█[0m[38;2;207;200;192m█[0m[38;2;202;197;191m█[0m[38;2;197;192;186m█[0m[38;2;193;186;180m█[0m[38;2;192;183;178m█[0m[38;2;193;185;174m█[0m[38;2;189;179;169m█[0m[38;2;190;180;171m█[0m[38;2;189;182;166m█[0m[38;2;186;174;158m█[0m[38;2;187;174;158m█[0m[38;2;184;171;155m█[0m[38;2;190;172;158m█[0m[38;2;189;171;157m█[0m[38;2;186;168;154m█[0m[38;2;181;169;155m█[0m[38;2;175;166;149m█[0m[38;2;168;162;140m█[0m[38;2;170;162;141m█[0m[38;2;172;160;136m█[0m[38;2;172;156;131m█[0m[38;2;177;161;135m█[0m[38;2;165;149;123m█[0m[38;2;169;153;127m█[0m[38;2;169;152;126m█[0m[38;2;168;151;125m█[0m[38;2;169;151;127m█[0m[38;2;172;152;128m█[0m[38;2;175;154;125m█[0m[38;2;178;155;123m█[0m[38;2;171;148;116m█[0m[38;2;173;150;118m█[0m[38;2;172;148;122m█[0m[38;2;176;152;126m█[0m[38;2;175;151;125m█[0m[38;2;174;150;114m█[0m[38;2;172;148;112m█[0m[38;2;167;143;107m█[0m[38;2;173;150;119m█[0m[38;2;170;150;123m█[0m[38;2;136;118;94m█[0m[38;2;0;0;0m██████[0m");
$display("[38;2;0;0;0m████████████████████████[0m[38;2;14;13;8m█[0m[38;2;117;116;98m█[0m[38;2;159;161;148m█[0m[38;2;138;132;136m█[0m[38;2;158;150;163m█[0m[38;2;216;208;219m█[0m[38;2;243;241;246m█[0m[38;2;240;242;241m█[0m[38;2;241;241;241m██[0m[38;2;240;240;240m█[0m[38;2;236;236;236m█[0m[38;2;230;232;231m█[0m[38;2;234;225;228m█[0m[38;2;228;222;224m█[0m[38;2;223;221;222m█[0m[38;2;227;218;221m█[0m[38;2;224;218;220m█[0m[38;2;226;222;223m█[0m[38;2;217;217;217m█[0m[38;2;221;221;221m█[0m[38;2;225;223;224m█[0m[38;2;228;222;224m█[0m[38;2;224;218;220m█[0m[38;2;218;213;209m█[0m[38;2;206;201;195m█[0m[38;2;196;191;185m█[0m[38;2;194;195;187m█[0m[38;2;195;190;184m█[0m[38;2;193;186;180m█[0m[38;2;191;186;180m█[0m[38;2;192;187;181m█[0m[38;2;189;186;179m█[0m[38;2;190;176;167m█[0m[38;2;185;175;165m█[0m[38;2;184;177;167m█[0m[38;2;184;175;168m█[0m[38;2;187;175;163m█[0m[38;2;188;174;161m█[0m[38;2;189;176;160m█[0m[38;2;184;171;155m███[0m[38;2;183;170;154m█[0m[38;2;182;169;153m█[0m[38;2;179;166;150m██[0m[38;2;178;165;149m█[0m[38;2;174;161;142m█[0m[38;2;168;156;130m█[0m[38;2;170;159;131m█[0m[38;2;175;158;132m█[0m[38;2;173;153;129m█[0m[38;2;171;152;135m█[0m[38;2;171;153;129m█[0m[38;2;172;155;129m█[0m[38;2;175;155;130m█[0m[38;2;174;152;128m█[0m[38;2;172;148;124m█[0m[38;2;175;151;127m█[0m[38;2;173;149;125m█[0m[38;2;168;143;121m█[0m[38;2;172;147;125m█[0m[38;2;173;148;126m█[0m[38;2;174;149;119m█[0m[38;2;172;147;117m█[0m[38;2;168;143;112m█[0m[38;2;167;147;120m█[0m[38;2;165;149;123m█[0m[38;2;134;119;96m█[0m[38;2;0;0;0m██████[0m");
$display("[38;2;0;0;0m████████████████████████[0m[38;2;29;30;25m█[0m[38;2;163;163;153m█[0m[38;2;146;155;154m█[0m[38;2;148;144;145m█[0m[38;2;198;189;194m█[0m[38;2;219;219;227m█[0m[38;2;240;239;244m█[0m[38;2;241;241;241m███[0m[38;2;239;239;239m█[0m[38;2;235;233;234m█[0m[38;2;231;227;228m█[0m[38;2;226;219;227m█[0m[38;2;213;207;209m█[0m[38;2;220;214;214m█[0m[38;2;215;209;209m█[0m[38;2;215;206;207m█[0m[38;2;216;207;208m█[0m[38;2;215;206;211m█[0m[38;2;214;212;215m█[0m[38;2;217;215;218m█[0m[38;2;222;222;224m█[0m[38;2;217;217;219m█[0m[38;2;208;204;201m█[0m[38;2;200;197;190m█[0m[38;2;194;192;180m█[0m[38;2;191;182;177m█[0m[38;2;188;179;170m█[0m[38;2;183;176;160m█[0m[38;2;183;175;164m███[0m[38;2;185;177;164m█[0m[38;2;186;178;165m█[0m[38;2;186;179;163m█[0m[38;2;185;178;160m█[0m[38;2;178;172;150m█[0m[38;2;182;174;153m█[0m[38;2;189;176;160m█[0m[38;2;186;173;157m█[0m[38;2;180;168;154m█[0m[38;2;181;173;154m█[0m[38;2;180;173;144m█[0m[38;2;179;170;153m█[0m[38;2;179;167;151m█[0m[38;2;178;169;152m█[0m[38;2;178;165;146m██[0m[38;2;171;160;138m█[0m[38;2;175;159;136m█[0m[38;2;180;158;137m█[0m[38;2;174;151;133m█[0m[38;2;174;155;140m█[0m[38;2;176;157;140m█[0m[38;2;175;157;137m█[0m[38;2;172;154;132m█[0m[38;2;170;146;122m█[0m[38;2;174;150;126m█[0m[38;2;172;148;120m█[0m[38;2;172;149;117m█[0m[38;2;170;145;115m█[0m[38;2;172;149;118m█[0m[38;2;168;149;117m█[0m[38;2;164;140;112m█[0m[38;2;166;142;116m█[0m[38;2;171;146;124m█[0m[38;2;170;155;126m█[0m[38;2;129;118;98m█[0m[38;2;0;0;0m███████[0m");
$display("[38;2;0;0;0m███████████████████████[0m[38;2;0;1;0m█[0m[38;2;195;189;191m█[0m[38;2;157;153;167m█[0m[38;2;125;121;135m█[0m[38;2;165;165;177m█[0m[38;2;212;212;224m█[0m[38;2;242;241;249m█[0m[38;2;243;243;245m█[0m[38;2;241;241;241m███[0m[38;2;236;236;236m█[0m[38;2;231;229;230m█[0m[38;2;231;222;225m█[0m[38;2;219;213;213m█[0m[38;2;211;206;203m█[0m[38;2;209;205;194m█[0m[38;2;203;199;188m█[0m[38;2;212;208;199m█[0m[38;2;210;206;197m█[0m[38;2;212;204;201m█[0m[38;2;207;206;201m█[0m[38;2;206;207;201m█[0m[38;2;217;216;211m█[0m[38;2;209;208;203m█[0m[38;2;197;194;189m█[0m[38;2;194;191;184m█[0m[38;2;181;182;168m█[0m[38;2;184;180;155m█[0m[38;2;180;173;154m█[0m[38;2;176;168;155m█[0m[38;2;171;162;153m█[0m[38;2;174;166;155m█[0m[38;2;181;172;163m█[0m[38;2;182;172;170m█[0m[38;2;182;173;168m██[0m[38;2;182;173;166m█[0m[38;2;179;171;158m█[0m[38;2;181;169;153m█[0m[38;2;186;170;155m█[0m[38;2;187;174;158m█[0m[38;2;182;173;158m████[0m[38;2;177;168;151m█[0m[38;2;174;167;149m█[0m[38;2;175;162;143m█[0m[38;2;177;164;145m█[0m[38;2;176;161;140m█[0m[38;2;177;158;143m█[0m[38;2;179;156;140m█[0m[38;2;182;156;141m█[0m[38;2;174;155;138m█[0m[38;2;175;156;139m█[0m[38;2;172;153;136m█[0m[38;2;176;155;134m█[0m[38;2;175;154;127m█[0m[38;2;175;151;127m█[0m[38;2;175;151;123m█[0m[38;2;172;152;119m█[0m[38;2;177;148;118m█[0m[38;2;169;148;117m█[0m[38;2;162;146;112m█[0m[38;2;163;139;111m█[0m[38;2;170;146;122m█[0m[38;2;173;151;128m█[0m[38;2;171;154;126m█[0m[38;2;156;141;118m█[0m[38;2;0;0;0m███████[0m");
$display("[38;2;0;0;0m███████████████████████[0m[38;2;4;4;4m█[0m[38;2;224;217;225m█[0m[38;2;184;181;192m█[0m[38;2;148;147;153m█[0m[38;2;191;190;196m█[0m[38;2;237;236;242m█[0m[38;2;241;241;241m██[0m[38;2;242;242;242m█[0m[38;2;243;243;243m█[0m[38;2;240;240;240m█[0m[38;2;230;230;230m█[0m[38;2;227;227;225m█[0m[38;2;214;215;209m█[0m[38;2;213;208;202m█[0m[38;2;197;192;186m█[0m[38;2;198;193;187m█[0m[38;2;199;194;188m█[0m[38;2;207;202;196m█[0m[38;2;209;204;198m█[0m[38;2;205;200;194m█[0m[38;2;207;202;196m█[0m[38;2;215;210;204m█[0m[38;2;212;207;201m█[0m[38;2;200;195;189m█[0m[38;2;188;183;177m█[0m[38;2;185;183;171m█[0m[38;2;176;173;158m█[0m[38;2;177;167;157m█[0m[38;2;173;165;154m█[0m[38;2;174;166;155m█[0m[38;2;174;165;158m█[0m[38;2;178;169;160m█[0m[38;2;176;167;160m█[0m[38;2;181;166;163m█[0m[38;2;182;172;163m█[0m[38;2;180;174;158m█[0m[38;2;179;172;153m█[0m[38;2;180;173;154m██[0m[38;2;182;170;154m█[0m[38;2;185;169;154m█[0m[38;2;187;169;155m█[0m[38;2;183;167;152m█[0m[38;2;182;164;150m█[0m[38;2;180;168;154m█[0m[38;2;176;163;146m█[0m[38;2;176;164;142m█[0m[38;2;176;163;146m█[0m[38;2;171;158;139m█[0m[38;2;169;157;135m█[0m[38;2;168;157;129m█[0m[38;2;173;155;135m█[0m[38;2;170;152;130m█[0m[38;2;169;151;127m█[0m[38;2;168;150;126m██[0m[38;2;167;149;125m█[0m[38;2;171;149;126m█[0m[38;2;173;149;125m█[0m[38;2;176;152;124m█[0m[38;2;172;149;117m█[0m[38;2;171;148;116m█[0m[38;2;168;144;118m█[0m[38;2;161;137;113m█[0m[38;2;162;134;113m█[0m[38;2;161;140;109m█[0m[38;2;164;146;124m█[0m[38;2;144;128;103m█[0m[38;2;74;66;55m█[0m[38;2;0;0;0m███████[0m");
$display("[38;2;0;0;0m██████████████████████[0m[38;2;1;1;1m█[0m[38;2;165;165;167m█[0m[38;2;207;212;216m█[0m[38;2;167;164;175m█[0m[38;2;161;160;168m█[0m[38;2;192;191;196m█[0m[38;2;240;240;242m█[0m[38;2;241;241;241m██[0m[38;2;244;244;244m█[0m[38;2;240;240;240m█[0m[38;2;235;235;235m█[0m[38;2;230;230;230m█[0m[38;2;216;216;214m█[0m[38;2;212;213;207m█[0m[38;2;208;203;197m█[0m[38;2;199;194;188m█[0m[38;2;193;188;182m█[0m[38;2;190;186;177m█[0m[38;2;191;187;176m█[0m[38;2;199;195;184m█[0m[38;2;196;196;188m██[0m[38;2;202;199;194m█[0m[38;2;201;196;192m█[0m[38;2;184;180;171m█[0m[38;2;183;181;168m█[0m[38;2;175;171;159m█[0m[38;2;175;165;155m█[0m[38;2;173;165;154m█[0m[38;2;171;163;152m█[0m[38;2;179;171;160m█[0m[38;2;176;170;154m█[0m[38;2;175;167;154m█[0m[38;2;179;165;152m█[0m[38;2;173;165;152m█[0m[38;2;169;162;146m█[0m[38;2;175;168;152m█[0m[38;2;178;171;155m█[0m[38;2;176;168;157m█[0m[38;2;181;173;162m█[0m[38;2;177;168;151m█[0m[38;2;182;173;156m█[0m[38;2;175;168;150m█[0m[38;2;171;162;145m█[0m[38;2;175;163;147m█[0m[38;2;179;163;150m█[0m[38;2;180;162;150m█[0m[38;2;179;163;148m█[0m[38;2;170;156;145m█[0m[38;2;173;156;136m█[0m[38;2;169;152;126m█[0m[38;2;169;158;130m█[0m[38;2;169;157;131m█[0m[38;2;160;145;122m█[0m[38;2;169;151;131m█[0m[38;2;168;150;130m█[0m[38;2;173;150;132m█[0m[38;2;171;146;126m█[0m[38;2;172;145;124m█[0m[38;2;174;150;126m█[0m[38;2;173;149;125m█[0m[38;2;171;147;119m█[0m[38;2;168;144;120m█[0m[38;2;163;136;115m█[0m[38;2;165;134;114m█[0m[38;2;167;140;113m█[0m[38;2;166;143;112m█[0m[38;2;170;149;130m█[0m[38;2;10;9;7m█[0m[38;2;0;0;0m████████[0m");
$display("[38;2;0;0;0m███████████████████████[0m[38;2;215;216;218m█[0m[38;2;231;238;244m█[0m[38;2;196;194;207m█[0m[38;2;165;164;172m█[0m[38;2;193;192;197m█[0m[38;2;237;237;239m█[0m[38;2;239;239;239m█[0m[38;2;241;241;241m█[0m[38;2;239;239;241m█[0m[38;2;234;234;234m█[0m[38;2;229;229;229m█[0m[38;2;227;227;229m█[0m[38;2;220;220;218m█[0m[38;2;212;213;207m█[0m[38;2;208;203;197m█[0m[38;2;197;192;186m█[0m[38;2;192;185;179m█[0m[38;2;191;185;173m█[0m[38;2;181;177;166m█[0m[38;2;185;178;170m█[0m[38;2;194;187;181m█[0m[38;2;188;179;174m█[0m[38;2;181;176;170m█[0m[38;2;180;174;162m█[0m[38;2;177;171;155m█[0m[38;2;172;170;155m█[0m[38;2;166;164;151m█[0m[38;2;164;156;145m█[0m[38;2;169;161;150m██[0m[38;2;172;164;153m█[0m[38;2;168;162;146m█[0m[38;2;170;158;144m█[0m[38;2;173;161;149m█[0m[38;2;176;169;153m█[0m[38;2;180;172;159m█[0m[38;2;177;170;152m█[0m[38;2;174;168;144m█[0m[38;2;178;171;153m█[0m[38;2;176;169;151m█[0m[38;2;177;165;149m█[0m[38;2;178;166;150m█[0m[38;2;174;167;149m█[0m[38;2;172;163;146m█[0m[38;2;177;165;149m█[0m[38;2;175;163;141m█[0m[38;2;159;149;124m█[0m[38;2;164;152;128m█[0m[38;2;160;154;130m█[0m[38;2;164;151;132m█[0m[38;2;163;150;133m█[0m[38;2;169;153;137m█[0m[38;2;162;149;132m█[0m[38;2;157;146;126m█[0m[38;2;160;147;128m██[0m[38;2;159;144;125m█[0m[38;2;161;143;121m█[0m[38;2;162;145;119m█[0m[38;2;164;142;118m█[0m[38;2;171;147;123m█[0m[38;2;171;147;121m█[0m[38;2;162;144;124m█[0m[38;2;161;139;118m█[0m[38;2;165;136;118m█[0m[38;2;161;141;117m█[0m[38;2;157;141;115m█[0m[38;2;95;86;79m█[0m[38;2;0;0;0m█████████[0m");
$display("[38;2;0;0;0m██████████████████████[0m[38;2;60;60;60m█[0m[38;2;235;234;240m█[0m[38;2;244;243;249m█[0m[38;2;202;201;207m█[0m[38;2;160;159;167m█[0m[38;2;222;221;226m█[0m[38;2;246;246;248m█[0m[38;2;242;241;246m█[0m[38;2;238;237;243m█[0m[38;2;234;233;239m█[0m[38;2;231;230;236m█[0m[38;2;233;232;238m█[0m[38;2;220;219;224m█[0m[38;2;215;215;215m█[0m[38;2;211;212;207m█[0m[38;2;199;199;191m█[0m[38;2;195;191;182m█[0m[38;2;196;188;175m█[0m[38;2;193;185;174m█[0m[38;2;184;176;165m█[0m[38;2;186;178;167m█[0m[38;2;182;174;163m█[0m[38;2;185;177;166m█[0m[38;2;182;174;163m█[0m[38;2;177;169;158m█[0m[38;2;171;163;152m█[0m[38;2;166;158;147m█[0m[38;2;168;160;149m█[0m[38;2;171;163;152m█[0m[38;2;168;161;142m█[0m[38;2;169;162;143m█[0m[38;2;165;158;139m█[0m[38;2;167;159;148m█[0m[38;2;168;160;149m█[0m[38;2;172;164;153m█[0m[38;2;171;162;157m█[0m[38;2;168;159;150m█[0m[38;2;172;165;149m█[0m[38;2;171;162;145m█[0m[38;2;165;156;139m█[0m[38;2;162;153;136m█[0m[38;2;169;156;140m█[0m[38;2;168;155;139m█[0m[38;2;168;156;140m█[0m[38;2;163;154;137m█[0m[38;2;164;155;138m█[0m[38;2;161;148;132m█[0m[38;2;170;157;141m█[0m[38;2;167;154;138m█[0m[38;2;166;153;134m█[0m[38;2;165;152;133m█[0m[38;2;147;136;116m█[0m[38;2;152;139;120m█[0m[38;2;157;140;122m█[0m[38;2;160;145;124m█[0m[38;2;155;143;117m█[0m[38;2;151;135;110m█[0m[38;2;151;133;111m█[0m[38;2;164;146;126m█[0m[38;2;163;145;121m█[0m[38;2;169;146;115m█[0m[38;2;168;145;114m█[0m[38;2;167;144;113m█[0m[38;2;164;137;118m█[0m[38;2;164;139;117m█[0m[38;2;155;137;113m█[0m[38;2;162;139;121m█[0m[38;2;154;141;122m█[0m[38;2;1;0;0m█[0m[38;2;0;0;0m█████████[0m");
$display("[38;2;0;0;0m██████████████████████[0m[38;2;161;161;163m█[0m[38;2;242;241;247m█[0m[38;2;238;237;243m█[0m[38;2;219;218;226m█[0m[38;2;173;172;180m█[0m[38;2;179;178;183m█[0m[38;2;231;231;233m█[0m[38;2;237;235;246m█[0m[38;2;234;233;241m█[0m[38;2;232;231;237m█[0m[38;2;229;228;234m█[0m[38;2;221;220;226m█[0m[38;2;217;218;213m█[0m[38;2;213;212;207m█[0m[38;2;212;208;197m█[0m[38;2;194;194;182m█[0m[38;2;194;190;179m█[0m[38;2;197;189;176m█[0m[38;2;198;190;177m█[0m[38;2;193;185;172m█[0m[38;2;188;180;167m█[0m[38;2;191;181;169m█[0m[38;2;187;177;165m█[0m[38;2;176;166;154m█[0m[38;2;171;161;151m██[0m[38;2;175;165;155m██[0m[38;2;172;162;152m█[0m[38;2;173;163;153m█[0m[38;2;171;161;152m█[0m[38;2;168;158;149m█[0m[38;2;164;155;150m█[0m[38;2;166;157;152m█[0m[38;2;169;160;153m█[0m[38;2;165;156;147m█[0m[38;2;161;154;144m█[0m[38;2;164;151;142m█[0m[38;2;165;155;146m█[0m[38;2;164;154;144m█[0m[38;2;160;150;138m█[0m[38;2;164;150;137m█[0m[38;2;164;148;135m█[0m[38;2;162;148;135m█[0m[38;2;167;149;135m█[0m[38;2;169;152;136m█[0m[38;2;164;152;136m█[0m[38;2;156;144;128m█[0m[38;2;163;151;135m█[0m[38;2;164;153;135m█[0m[38;2;160;149;131m█[0m[38;2;155;144;126m█[0m[38;2;147;136;116m█[0m[38;2;159;146;129m█[0m[38;2;155;142;123m█[0m[38;2;160;150;123m█[0m[38;2;161;145;120m█[0m[38;2;155;139;114m█[0m[38;2;153;137;111m██[0m[38;2;159;138;109m█[0m[38;2;163;142;113m█[0m[38;2;158;137;108m█[0m[38;2;166;140;115m█[0m[38;2;169;150;118m█[0m[38;2;165;149;124m█[0m[38;2;161;146;125m█[0m[38;2;56;49;43m█[0m[38;2;0;0;0m██████████[0m");
$display("\n");
$display("                                   \033[31m\033[5m █████ █████ █████ █████ █████ \033[0m");
$display("                                   \033[31m\033[5m █     █   █ █   █ █   █ █   █ \033[0m");
$display("                                   \033[31m\033[5m █████ █████ █████ █   █ █████ \033[0m");
$display("                                   \033[31m\033[5m █     █  █  █  █  █   █ █  █  \033[0m");
$display("                                   \033[31m\033[5m █████ █   █ █   █ █████ █   █ \033[0m");
$display("\n");

end endtask


task display_pass; begin

$display("[38;2;0;0;0m████████████████████████████████████████████████████[0m[38;2;1;1;1m█[0m[38;2;40;31;26m█[0m[38;2;68;57;53m█[0m[38;2;59;48;44m█[0m[38;2;26;16;15m█[0m[38;2;2;2;2m█[0m[38;2;0;1;0m█[0m[38;2;0;0;0m██████████████████████████████████████[0m");
$display("[38;2;0;0;0m███████████████████████████████████████████████████[0m[38;2;2;0;1m█[0m[38;2;0;1;3m█[0m[38;2;70;53;45m█[0m[38;2;72;44;30m█[0m[38;2;88;53;31m█[0m[38;2;100;55;36m█[0m[38;2;100;65;37m█[0m[38;2;101;65;41m█[0m[38;2;125;90;68m█[0m[38;2;113;85;71m█[0m[38;2;5;4;0m█[0m[38;2;0;0;0m███████████████████████████████████[0m");
$display("[38;2;0;0;0m████████████████████████████████████████████████████[0m[38;2;1;1;1m█[0m[38;2;30;16;15m█[0m[38;2;83;51;40m█[0m[38;2;101;59;34m█[0m[38;2;116;75;47m█[0m[38;2;125;84;54m█[0m[38;2;122;78;51m█[0m[38;2;109;67;42m█[0m[38;2;98;59;26m█[0m[38;2;98;69;39m█[0m[38;2;125;106;89m█[0m[38;2;16;8;5m█[0m[38;2;2;1;0m█[0m[38;2;1;1;3m█[0m[38;2;0;0;0m███████████████████████████████[0m");
$display("[38;2;0;0;0m█████████████[0m[38;2;254;0;0m█[0m[38;2;253;1;0m█[0m[38;2;200;20;31m█[0m[38;2;0;0;0m██[0m[38;2;0;7;4m█[0m[38;2;254;0;0m█[0m[38;2;0;3;2m█[0m[38;2;0;0;0m█[0m[38;2;254;1;0m█[0m[38;2;254;0;2m█[0m[38;2;0;0;0m███[0m[38;2;254;0;3m█[0m[38;2;254;0;0m████[0m[38;2;243;1;0m█[0m[38;2;0;0;0m██[0m[38;2;254;0;0m██████[0m[38;2;253;0;0m█[0m[38;2;0;0;0m███████████[0m[38;2;6;1;0m█[0m[38;2;95;63;50m█[0m[38;2;107;65;43m█[0m[38;2;120;78;53m█[0m[38;2;136;95;67m█[0m[38;2;137;93;66m█[0m[38;2;139;95;68m█[0m[38;2;135;94;62m█[0m[38;2;115;77;41m█[0m[38;2;102;65;36m█[0m[38;2;98;71;44m█[0m[38;2;92;76;60m█[0m[38;2;0;0;0m█[0m[38;2;3;3;3m█[0m[38;2;0;0;0m██████████████████████████████[0m");
$display("[38;2;0;0;0m█████████████[0m[38;2;254;0;0m█[0m[38;2;254;0;5m█[0m[38;2;254;0;0m█[0m[38;2;245;3;1m█[0m[38;2;0;1;0m█[0m[38;2;0;7;4m█[0m[38;2;254;0;0m█[0m[38;2;0;3;2m█[0m[38;2;0;0;0m█[0m[38;2;254;1;0m█[0m[38;2;254;0;2m█[0m[38;2;0;0;0m█[0m[38;2;1;0;0m█[0m[38;2;254;0;0m█[0m[38;2;254;2;0m█[0m[38;2;0;0;0m███[0m[38;2;18;0;0m█[0m[38;2;0;0;0m███[0m[38;2;254;0;0m██[0m[38;2;3;0;0m████[0m[38;2;0;0;0m████████████[0m[38;2;2;1;7m█[0m[38;2;58;39;25m█[0m[38;2;104;64;39m█[0m[38;2;121;77;50m█[0m[38;2;127;83;54m█[0m[38;2;131;89;64m█[0m[38;2;139;102;75m█[0m[38;2;145;108;79m█[0m[38;2;143;106;77m█[0m[38;2;137;101;69m█[0m[38;2;112;73;40m█[0m[38;2;99;65;38m█[0m[38;2;111;84;63m█[0m[38;2;56;48;37m█[0m[38;2;0;2;1m█[0m[38;2;1;1;1m█[0m[38;2;0;0;0m████████████████████████████[0m");
$display("[38;2;0;0;0m█████████████[0m[38;2;254;0;0m█[0m[38;2;254;0;2m█[0m[38;2;6;0;0m█[0m[38;2;248;2;5m█[0m[38;2;254;0;0m█[0m[38;2;0;6;4m█[0m[38;2;254;0;0m█[0m[38;2;0;3;2m█[0m[38;2;0;0;0m█[0m[38;2;254;1;0m█[0m[38;2;254;0;2m█[0m[38;2;0;0;0m█[0m[38;2;166;22;21m█[0m[38;2;254;0;0m█[0m[38;2;0;0;0m████████[0m[38;2;254;0;0m██[0m[38;2;254;0;2m████[0m[38;2;0;0;0m████████████[0m[38;2;1;1;1m██[0m[38;2;78;49;35m█[0m[38;2;129;85;58m█[0m[38;2;150;101;71m█[0m[38;2;145;100;71m█[0m[38;2;152;113;84m█[0m[38;2;150;115;83m█[0m[38;2;145;112;79m█[0m[38;2;142;107;75m█[0m[38;2;140;105;75m█[0m[38;2;134;98;72m█[0m[38;2;109;73;47m█[0m[38;2;110;77;46m█[0m[38;2;109;88;67m█[0m[38;2;60;51;46m█[0m[38;2;0;0;4m█[0m[38;2;0;0;0m█[0m[38;2;0;0;2m█[0m[38;2;0;0;0m█████████████████████████[0m");
$display("[38;2;0;0;0m█████████████[0m[38;2;254;0;0m██[0m[38;2;0;0;0m█[0m[38;2;0;0;4m█[0m[38;2;247;3;2m█[0m[38;2;254;0;0m██[0m[38;2;0;3;2m█[0m[38;2;0;0;0m█[0m[38;2;254;1;0m█[0m[38;2;254;0;2m█[0m[38;2;0;0;0m█[0m[38;2;9;0;0m█[0m[38;2;251;1;2m█[0m[38;2;251;0;0m█[0m[38;2;0;0;0m███[0m[38;2;250;0;3m█[0m[38;2;254;0;2m█[0m[38;2;11;1;2m█[0m[38;2;0;0;0m█[0m[38;2;254;0;0m██[0m[38;2;0;0;0m██████████████████[0m[38;2;34;17;7m█[0m[38;2;86;60;37m█[0m[38;2;125;87;64m█[0m[38;2;133;92;60m█[0m[38;2;138;103;75m█[0m[38;2;145;113;90m█[0m[38;2;152;115;88m█[0m[38;2;148;112;86m█[0m[38;2;152;116;90m█[0m[38;2;147;111;85m█[0m[38;2;142;106;82m█[0m[38;2;133;94;61m█[0m[38;2;93;58;38m█[0m[38;2;109;78;58m█[0m[38;2;126;98;84m█[0m[38;2;85;65;56m█[0m[38;2;7;2;0m█[0m[38;2;2;1;0m█[0m[38;2;7;7;5m█[0m[38;2;11;9;10m██[0m[38;2;9;7;8m█[0m[38;2;11;9;10m█[0m[38;2;28;22;22m█[0m[38;2;36;32;31m█[0m[38;2;65;60;64m█[0m[38;2;77;74;67m█[0m[38;2;66;63;58m█[0m[38;2;50;47;40m█[0m[38;2;40;37;32m█[0m[38;2;49;45;42m█[0m[38;2;41;37;36m█[0m[38;2;12;10;11m█[0m[38;2;1;1;0m█[0m[38;2;0;0;2m█[0m[38;2;1;1;1m█[0m[38;2;0;0;4m█[0m[38;2;1;1;1m██[0m[38;2;1;1;3m██[0m[38;2;78;73;69m█[0m");
$display("[38;2;0;0;0m█████████████[0m[38;2;254;0;0m██[0m[38;2;0;0;0m███[0m[38;2;254;0;0m██[0m[38;2;0;3;2m█[0m[38;2;0;0;0m█[0m[38;2;254;1;0m█[0m[38;2;254;0;2m█[0m[38;2;0;0;0m██[0m[38;2;6;0;0m█[0m[38;2;254;0;0m██[0m[38;2;253;1;0m█[0m[38;2;254;0;0m██[0m[38;2;0;5;4m█[0m[38;2;0;0;0m██[0m[38;2;254;0;0m██████[0m[38;2;254;0;7m█[0m[38;2;0;0;0m█████████████[0m[38;2;32;25;19m█[0m[38;2;123;108;87m█[0m[38;2;141;115;90m█[0m[38;2;157;124;93m█[0m[38;2;153;121;96m█[0m[38;2;152;125;96m█[0m[38;2;160;133;104m█[0m[38;2;161;130;102m█[0m[38;2;159;128;100m█[0m[38;2;161;130;102m█[0m[38;2;148;116;91m█[0m[38;2;134;102;79m█[0m[38;2;98;66;45m█[0m[38;2;101;69;48m█[0m[38;2;126;91;71m█[0m[38;2;104;83;56m█[0m[38;2;48;33;4m█[0m[38;2;67;49;27m█[0m[38;2;61;41;30m█[0m[38;2;51;34;27m█[0m[38;2;36;20;20m█[0m[38;2;29;19;18m█[0m[38;2;31;21;22m█[0m[38;2;27;17;18m██[0m[38;2;31;21;22m█[0m[38;2;24;14;15m█[0m[38;2;28;18;19m█[0m[38;2;40;30;31m█[0m[38;2;29;21;18m█[0m[38;2;20;16;7m█[0m[38;2;33;29;17m█[0m[38;2;39;27;15m█[0m[38;2;49;35;22m█[0m[38;2;52;45;26m█[0m[38;2;70;59;39m█[0m[38;2;87;61;46m█[0m[38;2;106;78;64m█[0m[38;2;116;87;73m█[0m[38;2;128;105;87m█[0m[38;2;107;85;71m█[0m[38;2;78;57;40m█[0m");
$display("[38;2;0;0;0m███████████████████████████████████████████████████████[0m[38;2;5;0;0m█[0m[38;2;115;107;86m█[0m[38;2;139;111;87m█[0m[38;2;184;149;119m█[0m[38;2;181;150;122m█[0m[38;2;171;146;116m█[0m[38;2;164;139;109m█[0m[38;2;163;137;110m█[0m[38;2;163;135;111m█[0m[38;2;163;133;107m█[0m[38;2;153;122;94m█[0m[38;2;145;110;91m█[0m[38;2;123;91;70m█[0m[38;2;118;90;66m█[0m[38;2;98;77;46m█[0m[38;2;100;83;55m█[0m[38;2;78;67;39m█[0m[38;2;51;41;16m█[0m[38;2;43;31;15m█[0m[38;2;34;22;8m█[0m[38;2;38;29;20m█[0m[38;2;32;22;21m█[0m[38;2;40;29;33m█[0m[38;2;33;22;26m█[0m[38;2;32;22;21m█[0m[38;2;48;38;39m█[0m[38;2;46;35;41m█[0m[38;2;45;35;34m█[0m[38;2;54;44;43m█[0m[38;2;20;12;9m█[0m[38;2;33;29;20m█[0m[38;2;39;36;29m█[0m[38;2;29;31;17m█[0m[38;2;38;35;18m█[0m[38;2;56;50;28m█[0m[38;2;42;29;13m█[0m[38;2;50;27;13m█[0m[38;2;77;50;31m█[0m[38;2;119;92;73m█[0m[38;2;96;67;53m█[0m[38;2;74;45;31m█[0m[38;2;86;57;43m█[0m");
$display("[38;2;0;0;0m███████████████████████████████████████████████████████[0m[38;2;3;1;2m█[0m[38;2;140;135;113m█[0m[38;2;166;142;114m█[0m[38;2;178;138;112m█[0m[38;2;185;147;126m█[0m[38;2;171;140;111m█[0m[38;2;157;132;101m█[0m[38;2;156;131;101m█[0m[38;2;158;133;103m█[0m[38;2;160;135;105m█[0m[38;2;150;125;94m█[0m[38;2;142;115;88m█[0m[38;2;137;106;77m█[0m[38;2;111;84;54m█[0m[38;2;86;62;36m█[0m[38;2;68;53;32m█[0m[38;2;36;26;14m█[0m[38;2;25;17;4m█[0m[38;2;31;24;8m█[0m[38;2;48;41;31m█[0m[38;2;43;39;30m█[0m[38;2;48;39;34m█[0m[38;2;82;73;68m█[0m[38;2;50;41;34m█[0m[38;2;19;11;0m█[0m[38;2;46;37;28m█[0m[38;2;46;37;30m█[0m[38;2;41;32;25m█[0m[38;2;40;31;24m█[0m[38;2;35;25;16m█[0m[38;2;34;24;14m█[0m[38;2;42;39;24m█[0m[38;2;50;41;24m█[0m[38;2;64;51;34m█[0m[38;2;58;42;17m█[0m[38;2;84;66;42m█[0m[38;2;128;100;79m█[0m[38;2;113;81;60m█[0m[38;2;108;76;55m█[0m[38;2;93;58;36m█[0m[38;2;101;66;44m█[0m[38;2;106;71;49m█[0m");
$display("[38;2;0;0;0m███████████████████████████████████████████████████████[0m[38;2;4;0;0m█[0m[38;2;121;104;86m█[0m[38;2;139;104;85m█[0m[38;2;174;126;103m█[0m[38;2;178;134;109m█[0m[38;2;178;139;108m█[0m[38;2;166;136;102m█[0m[38;2;151;120;89m█[0m[38;2;147;118;88m█[0m[38;2;157;132;102m█[0m[38;2;141;118;87m█[0m[38;2;134;108;75m█[0m[38;2;121;95;72m█[0m[38;2;87;63;39m█[0m[38;2;67;49;25m█[0m[38;2;51;34;14m█[0m[38;2;23;20;1m█[0m[38;2;33;24;7m█[0m[38;2;64;55;38m█[0m[38;2;89;81;68m█[0m[38;2;105;97;84m█[0m[38;2;100;91;82m█[0m[38;2;101;92;83m█[0m[38;2;64;55;46m█[0m[38;2;60;52;41m█[0m[38;2;53;44;35m█[0m[38;2;48;39;30m█[0m[38;2;39;35;24m█[0m[38;2;28;24;13m█[0m[38;2;27;18;9m█[0m[38;2;55;38;30m█[0m[38;2;78;55;47m█[0m[38;2;81;55;40m█[0m[38;2;74;51;35m█[0m[38;2;94;68;43m█[0m[38;2;110;82;60m█[0m[38;2;133;96;77m█[0m[38;2;131;91;65m█[0m[38;2;134;94;68m█[0m[38;2;138;102;70m█[0m[38;2;134;102;77m█[0m[38;2;115;83;62m█[0m");
$display("[38;2;0;0;0m█████[0m[38;2;2;0;3m█[0m[38;2;254;1;0m██[0m[38;2;254;0;0m█[0m[38;2;254;0;2m█[0m[38;2;254;1;0m█[0m[38;2;249;0;0m█[0m[38;2;0;4;0m█[0m[38;2;0;0;0m█[0m[38;2;0;8;2m█[0m[38;2;254;0;0m█[0m[38;2;249;7;0m█[0m[38;2;0;0;0m███[0m[38;2;254;1;0m█[0m[38;2;254;0;0m█[0m[38;2;10;0;0m█[0m[38;2;0;7;0m█[0m[38;2;254;1;0m██[0m[38;2;254;0;0m██[0m[38;2;250;3;0m█[0m[38;2;225;14;21m█[0m[38;2;0;0;2m█[0m[38;2;0;0;0m██[0m[38;2;254;1;0m██[0m[38;2;254;0;0m██[0m[38;2;251;3;0m█[0m[38;2;255;5;0m█[0m[38;2;4;0;0m█[0m[38;2;0;0;0m█[0m[38;2;13;0;0m█[0m[38;2;254;1;0m█[0m[38;2;254;2;0m█[0m[38;2;0;1;2m█[0m[38;2;0;0;0m██[0m[38;2;8;0;2m█[0m[38;2;254;0;0m█[0m[38;2;251;0;0m█[0m[38;2;0;4;0m█[0m[38;2;0;0;0m████[0m[38;2;2;1;0m█[0m[38;2;153;131;117m█[0m[38;2;159;120;105m█[0m[38;2;161;113;93m█[0m[38;2;158;117;89m█[0m[38;2;143;107;75m█[0m[38;2;143;110;77m█[0m[38;2;138;107;76m█[0m[38;2;134;103;74m█[0m[38;2;122;92;64m█[0m[38;2;93;68;38m█[0m[38;2;99;74;44m█[0m[38;2;90;66;42m█[0m[38;2;85;59;34m█[0m[38;2;110;80;52m█[0m[38;2;109;88;67m█[0m[38;2;95;82;65m█[0m[38;2;127;120;102m█[0m[38;2;158;151;133m█[0m[38;2;139;130;115m█[0m[38;2;183;174;159m█[0m[38;2;181;173;162m█[0m[38;2;144;136;123m█[0m[38;2;140;132;119m█[0m[38;2;120;112;99m█[0m[38;2;61;53;40m█[0m[38;2;30;22;9m█[0m[38;2;48;42;28m█[0m[38;2;67;61;47m█[0m[38;2;59;49;37m█[0m[38;2;69;52;42m█[0m[38;2;59;35;23m█[0m[38;2;47;21;8m█[0m[38;2;88;62;47m█[0m[38;2;81;56;34m█[0m[38;2;96;68;46m█[0m[38;2;104;68;44m█[0m[38;2;111;75;49m█[0m[38;2;147;111;85m█[0m[38;2;152;118;90m█[0m[38;2;144;113;85m█[0m[38;2;136;104;79m█[0m");
$display("[38;2;0;0;0m█████[0m[38;2;0;5;0m█[0m[38;2;254;0;0m█[0m[38;2;160;0;0m█[0m[38;2;0;0;2m█[0m[38;2;0;0;5m█[0m[38;2;0;3;2m█[0m[38;2;254;0;0m██[0m[38;2;0;0;0m█[0m[38;2;0;2;4m█[0m[38;2;254;0;0m█[0m[38;2;251;3;4m█[0m[38;2;0;0;0m███[0m[38;2;247;4;0m█[0m[38;2;254;0;0m█[0m[38;2;8;0;0m█[0m[38;2;0;1;2m█[0m[38;2;254;0;0m██[0m[38;2;0;1;0m█[0m[38;2;0;0;4m█[0m[38;2;0;0;0m█[0m[38;2;237;11;0m█[0m[38;2;254;0;0m█[0m[38;2;9;0;3m█[0m[38;2;0;0;0m█[0m[38;2;254;0;0m██[0m[38;2;1;0;0m█[0m[38;2;0;0;0m█[0m[38;2;0;0;4m█[0m[38;2;234;8;19m█[0m[38;2;254;0;0m█[0m[38;2;132;4;0m█[0m[38;2;0;0;0m█[0m[38;2;3;0;5m█[0m[38;2;254;0;0m█[0m[38;2;254;0;2m█[0m[38;2;0;2;0m█[0m[38;2;0;0;0m█[0m[38;2;254;0;0m█[0m[38;2;254;2;0m█[0m[38;2;0;0;0m████[0m[38;2;2;0;3m█[0m[38;2;0;0;0m█[0m[38;2;130;113;103m█[0m[38;2;179;153;136m█[0m[38;2;156;118;109m█[0m[38;2;157;111;88m█[0m[38;2;150;110;85m█[0m[38;2;131;95;69m█[0m[38;2;132;98;71m█[0m[38;2;131;95;69m█[0m[38;2;112;75;49m█[0m[38;2;132;97;77m█[0m[38;2;134;106;85m█[0m[38;2;120;102;82m█[0m[38;2;115;94;77m█[0m[38;2;114;96;74m█[0m[38;2;150;129;108m█[0m[38;2;145;129;106m█[0m[38;2;155;139;123m█[0m[38;2;191;178;162m█[0m[38;2;197;184;168m█[0m[38;2;192;185;167m█[0m[38;2;196;189;171m█[0m[38;2;199;192;174m█[0m[38;2;187;180;162m█[0m[38;2;180;173;155m█[0m[38;2;144;137;119m█[0m[38;2;91;82;65m█[0m[38;2;58;49;32m█[0m[38;2;87;74;58m█[0m[38;2;91;78;62m█[0m[38;2;103;85;71m█[0m[38;2;102;83;66m█[0m[38;2;87;64;46m█[0m[38;2;63;37;20m█[0m[38;2;72;46;31m█[0m[38;2;63;38;16m█[0m[38;2;78;51;30m█[0m[38;2;79;52;31m█[0m[38;2;89;58;30m█[0m[38;2;96;65;37m█[0m[38;2;102;75;46m█[0m[38;2;123;98;68m██[0m");
$display("[38;2;0;0;0m█████[0m[38;2;0;5;0m█[0m[38;2;254;0;0m█████[0m[38;2;255;5;3m█[0m[38;2;4;0;0m█[0m[38;2;0;0;0m█[0m[38;2;0;2;4m█[0m[38;2;254;0;0m█[0m[38;2;248;4;4m█[0m[38;2;0;0;0m███[0m[38;2;247;4;0m█[0m[38;2;254;0;0m█[0m[38;2;10;0;0m█[0m[38;2;0;1;2m█[0m[38;2;254;0;0m██[0m[38;2;0;2;2m█[0m[38;2;0;0;0m██[0m[38;2;14;0;0m█[0m[38;2;254;0;0m██[0m[38;2;0;0;0m█[0m[38;2;254;0;0m██[0m[38;2;4;0;0m█[0m[38;2;0;0;0m██[0m[38;2;1;0;5m█[0m[38;2;254;0;0m██[0m[38;2;0;0;0m███[0m[38;2;250;3;0m█[0m[38;2;254;0;0m█[0m[38;2;248;4;0m█[0m[38;2;171;7;8m█[0m[38;2;0;0;0m█████[0m[38;2;4;0;3m█[0m[38;2;4;0;1m█[0m[38;2;173;147;134m█[0m[38;2;175;145;121m█[0m[38;2;164;129;109m█[0m[38;2;147;109;86m█[0m[38;2;144;107;81m█[0m[38;2;122;88;61m█[0m[38;2;124;95;61m█[0m[38;2;124;97;68m█[0m[38;2;101;75;50m█[0m[38;2;109;85;61m█[0m[38;2;138;110;99m█[0m[38;2;117;98;84m█[0m[38;2;134;115;101m█[0m[38;2;149;131;117m█[0m[38;2;183;170;154m█[0m[38;2;189;177;161m█[0m[38;2;183;171;155m█[0m[38;2;188;179;162m█[0m[38;2;196;187;170m█[0m[38;2;197;188;171m█[0m[38;2;200;191;174m█[0m[38;2;197;188;171m█[0m[38;2;202;193;176m█[0m[38;2;198;189;172m█[0m[38;2;174;169;150m█[0m[38;2;173;166;148m█[0m[38;2;125;118;100m█[0m[38;2;97;88;71m█[0m[38;2;93;84;67m█[0m[38;2;105;100;81m█[0m[38;2;108;96;80m█[0m[38;2;103;80;66m█[0m[38;2;133;106;89m█[0m[38;2;114;86;72m█[0m[38;2;106;79;62m█[0m[38;2;93;66;49m█[0m[38;2;107;80;63m█[0m[38;2;98;74;48m█[0m[38;2;96;75;48m█[0m[38;2;98;72;47m█[0m[38;2;99;78;51m█[0m[38;2;94;77;49m█[0m");
$display("[38;2;0;0;0m█████[0m[38;2;0;5;0m█[0m[38;2;254;0;0m█[0m[38;2;158;0;0m█[0m[38;2;0;0;0m███[0m[38;2;251;3;0m█[0m[38;2;254;0;0m█[0m[38;2;0;0;0m█[0m[38;2;0;3;5m█[0m[38;2;254;0;0m█[0m[38;2;245;1;0m█[0m[38;2;0;0;0m███[0m[38;2;250;1;5m█[0m[38;2;254;0;0m█[0m[38;2;4;0;2m█[0m[38;2;0;1;2m█[0m[38;2;254;0;0m██[0m[38;2;0;2;2m█[0m[38;2;0;0;0m██[0m[38;2;0;6;7m█[0m[38;2;254;0;0m█[0m[38;2;254;0;2m█[0m[38;2;0;0;0m█[0m[38;2;254;0;0m██[0m[38;2;4;0;0m█[0m[38;2;0;0;0m██[0m[38;2;7;0;0m█[0m[38;2;254;0;0m██[0m[38;2;0;0;0m████[0m[38;2;251;2;0m█[0m[38;2;255;1;0m█[0m[38;2;0;0;0m██████[0m[38;2;1;1;1m██[0m[38;2;157;131;114m█[0m[38;2;165;131;106m█[0m[38;2;153;121;98m█[0m[38;2;142;110;85m█[0m[38;2;128;98;70m█[0m[38;2;126;97;67m█[0m[38;2;120;100;63m█[0m[38;2;125;102;70m█[0m[38;2;128;104;78m█[0m[38;2;172;147;125m█[0m[38;2;149;123;110m█[0m[38;2;146;127;113m█[0m[38;2;156;132;120m█[0m[38;2;186;168;154m█[0m[38;2;186;173;157m█[0m[38;2;185;172;156m██[0m[38;2;189;177;161m█[0m[38;2;191;179;163m█[0m[38;2;192;183;166m█[0m[38;2;196;184;168m█[0m[38;2;198;189;172m█[0m[38;2;200;188;172m█[0m[38;2;200;191;174m█[0m[38;2;205;198;180m█[0m[38;2;202;195;177m█[0m[38;2;147;140;122m█[0m[38;2;92;83;66m█[0m[38;2;120;111;94m█[0m[38;2;107;102;83m█[0m[38;2;108;91;75m█[0m[38;2;77;54;40m█[0m[38;2;89;62;45m█[0m[38;2;94;66;52m█[0m[38;2;65;37;23m█[0m[38;2;91;64;47m█[0m[38;2;100;73;56m█[0m[38;2;91;65;42m█[0m[38;2;94;68;45m█[0m[38;2;97;71;48m█[0m[38;2;105;79;56m█[0m[38;2;104;80;56m█[0m");
$display("[38;2;0;0;0m█████[0m[38;2;0;5;0m█[0m[38;2;254;0;0m█[0m[38;2;254;0;7m█[0m[38;2;240;7;3m█[0m[38;2;241;5;9m█[0m[38;2;254;3;0m█[0m[38;2;254;0;0m██[0m[38;2;0;0;0m█[0m[38;2;0;1;5m█[0m[38;2;253;0;0m█[0m[38;2;254;0;0m█[0m[38;2;254;1;0m█[0m[38;2;22;0;0m█[0m[38;2;254;1;0m█[0m[38;2;254;0;0m█[0m[38;2;247;5;0m█[0m[38;2;0;2;0m█[0m[38;2;0;1;2m█[0m[38;2;254;0;0m██[0m[38;2;240;7;3m█[0m[38;2;246;4;3m█[0m[38;2;254;1;0m█[0m[38;2;254;0;0m█[0m[38;2;245;0;0m█[0m[38;2;0;8;2m█[0m[38;2;0;0;0m█[0m[38;2;254;0;0m██[0m[38;2;237;7;9m█[0m[38;2;241;6;3m█[0m[38;2;254;1;0m█[0m[38;2;254;0;0m█[0m[38;2;251;0;0m█[0m[38;2;3;0;11m█[0m[38;2;0;0;0m████[0m[38;2;251;2;0m█[0m[38;2;254;1;0m█[0m[38;2;0;0;0m██████[0m[38;2;3;1;4m█[0m[38;2;84;67;57m█[0m[38;2;130;95;75m█[0m[38;2;126;92;64m█[0m[38;2;139;105;78m█[0m[38;2;136;107;77m█[0m[38;2;144;117;87m█[0m[38;2;145;120;89m█[0m[38;2;155;130;99m█[0m[38;2;144;118;93m█[0m[38;2;151;125;108m█[0m[38;2;180;157;143m█[0m[38;2;168;141;130m█[0m[38;2;160;142;128m█[0m[38;2;182;163;149m█[0m[38;2;182;164;150m█[0m[38;2;175;162;146m█[0m[38;2;182;169;153m█[0m[38;2;187;174;158m█[0m[38;2;188;176;160m█[0m[38;2;193;181;165m█[0m[38;2;198;186;170m█[0m[38;2;191;179;163m█[0m[38;2;203;190;174m█[0m[38;2;201;188;172m█[0m[38;2;200;188;172m█[0m[38;2;204;197;179m█[0m[38;2;206;197;180m█[0m[38;2;192;183;166m█[0m[38;2;133;124;107m█[0m[38;2;148;139;122m█[0m[38;2;144;137;118m█[0m[38;2;135;118;98m█[0m[38;2;111;88;72m█[0m[38;2;125;98;81m█[0m[38;2;122;94;80m█[0m[38;2;106;78;64m█[0m[38;2;101;73;59m█[0m[38;2;103;75;61m█[0m[38;2;109;83;60m█[0m[38;2;103;77;54m█[0m[38;2;98;72;49m█[0m[38;2;94;68;45m█[0m[38;2;97;71;48m█[0m");
$display("[38;2;0;0;0m█████[0m[38;2;6;0;0m█[0m[38;2;0;0;0m███[0m[38;2;3;0;2m█[0m[38;2;3;0;0m█[0m[38;2;0;3;4m█[0m[38;2;0;0;0m████[0m[38;2;0;2;5m█[0m[38;2;4;0;0m█[0m[38;2;18;0;0m█[0m[38;2;1;0;0m█[0m[38;2;3;0;0m█[0m[38;2;0;0;0m██[0m[38;2;1;0;2m█[0m[38;2;0;0;0m███[0m[38;2;0;2;0m█[0m[38;2;3;0;0m██[0m[38;2;0;0;0m██[0m[38;2;0;1;0m█[0m[38;2;0;0;0m████[0m[38;2;0;0;4m█[0m[38;2;6;0;0m█[0m[38;2;0;0;0m███████[0m[38;2;3;0;7m█[0m[38;2;0;0;0m████[0m[38;2;0;0;4m█[0m[38;2;12;11;6m█[0m[38;2;68;54;43m█[0m[38;2;105;88;68m█[0m[38;2;121;102;70m█[0m[38;2;118;97;70m█[0m[38;2;112;91;70m█[0m[38;2;111;96;77m█[0m[38;2;114;103;85m█[0m[38;2;118;106;80m█[0m[38;2;131;118;99m█[0m[38;2;123;112;92m█[0m[38;2;140;127;111m█[0m[38;2;149;130;116m█[0m[38;2;156;137;123m█[0m[38;2;168;150;136m█[0m[38;2;176;154;141m█[0m[38;2;179;160;146m█[0m[38;2;186;167;153m█[0m[38;2;189;170;156m██[0m[38;2;190;171;157m█[0m[38;2;198;179;165m█[0m[38;2;203;184;170m█[0m[38;2;199;180;166m█[0m[38;2;203;184;170m█[0m[38;2;209;190;176m█[0m[38;2;206;187;173m█[0m[38;2;204;188;173m█[0m[38;2;202;186;171m█[0m[38;2;203;190;174m█[0m[38;2;208;199;182m█[0m[38;2;185;176;159m█[0m[38;2;160;152;133m█[0m[38;2;148;133;114m█[0m[38;2;120;97;81m█[0m[38;2;126;98;84m█[0m[38;2;115;87;73m█[0m[38;2;101;73;59m█[0m[38;2;110;82;70m█[0m[38;2;114;86;74m█[0m[38;2;127;101;78m█[0m[38;2;124;98;75m█[0m[38;2;118;92;69m█[0m[38;2;114;88;65m█[0m[38;2;103;77;54m█[0m");
$display("[38;2;0;0;0m█████████████████████████████████████████████████[0m[38;2;1;1;1m█[0m[38;2;3;2;0m█[0m[38;2;49;35;22m█[0m[38;2;74;47;38m█[0m[38;2;81;64;54m█[0m[38;2;86;70;54m█[0m[38;2;84;72;48m█[0m[38;2;80;70;43m█[0m[38;2;61;48;39m█[0m[38;2;40;32;29m█[0m[38;2;35;30;27m█[0m[38;2;22;23;28m█[0m[38;2;26;27;22m█[0m[38;2;28;31;22m█[0m[38;2;90;92;78m█[0m[38;2;72;64;53m█[0m[38;2;109;92;84m█[0m[38;2;133;115;105m█[0m[38;2;163;144;130m█[0m[38;2;180;161;147m█[0m[38;2;182;163;149m█[0m[38;2;190;171;157m█[0m[38;2;188;169;155m█[0m[38;2;195;176;162m█[0m[38;2;201;182;168m█[0m[38;2;204;185;171m█[0m[38;2;203;184;170m█[0m[38;2;204;185;171m██[0m[38;2;198;180;166m█[0m[38;2;194;176;162m█[0m[38;2;202;180;167m█[0m[38;2;197;184;168m█[0m[38;2;182;173;156m█[0m[38;2;179;170;153m█[0m[38;2;162;147;128m█[0m[38;2;157;145;123m█[0m[38;2;145;128;108m█[0m[38;2;156;128;114m█[0m[38;2;158;130;118m█[0m[38;2;154;126;104m█[0m[38;2;142;110;89m█[0m[38;2;131;100;79m█[0m[38;2;111;79;58m█[0m[38;2;126;94;73m█[0m[38;2;118;90;68m█[0m[38;2;115;88;67m█[0m[38;2;114;87;66m█[0m");
$display("[38;2;0;0;0m█████████████████████████████████████████████████[0m[38;2;21;17;18m█[0m[38;2;101;86;79m█[0m[38;2;90;71;57m██[0m[38;2;95;79;64m█[0m[38;2;117;104;88m█[0m[38;2;120;107;88m█[0m[38;2;95;87;66m█[0m[38;2;44;35;26m█[0m[38;2;30;20;21m█[0m[38;2;25;20;27m█[0m[38;2;19;22;29m█[0m[38;2;20;24;35m█[0m[38;2;42;47;50m█[0m[38;2;39;44;38m█[0m[38;2;61;65;51m█[0m[38;2;57;50;40m█[0m[38;2;105;86;72m█[0m[38;2;144;124;113m█[0m[38;2;165;147;133m█[0m[38;2;178;160;146m█[0m[38;2;188;170;156m█[0m[38;2;197;173;161m█[0m[38;2;200;181;167m█[0m[38;2;198;179;165m█[0m[38;2;204;185;171m█[0m[38;2;202;183;169m█[0m[38;2;204;182;169m█[0m[38;2;206;184;171m██[0m[38;2;196;177;163m█[0m[38;2;190;170;159m█[0m[38;2;187;171;156m█[0m[38;2;176;164;148m█[0m[38;2;160;149;131m█[0m[38;2;148;135;116m█[0m[38;2;142;127;108m█[0m[38;2;136;125;105m█[0m[38;2;114;106;85m█[0m[38;2;84;69;50m█[0m[38;2;88;67;46m█[0m[38;2;127;103;79m█[0m[38;2;157;125;102m█[0m[38;2;153;122;101m█[0m[38;2;131;99;76m█[0m[38;2;112;82;58m█[0m[38;2;97;69;48m█[0m[38;2;116;90;67m█[0m");
$display("[38;2;0;0;0m████████████████████████████████████████████████[0m[38;2;9;3;3m█[0m[38;2;105;85;74m█[0m[38;2;93;69;57m█[0m[38;2;75;56;42m█[0m[38;2;76;57;43m█[0m[38;2;91;82;65m█[0m[38;2;122;113;96m█[0m[38;2;124;116;103m█[0m[38;2;89;86;71m█[0m[38;2;40;36;35m█[0m[38;2;15;13;18m█[0m[38;2;27;24;33m█[0m[38;2;32;32;42m█[0m[38;2;42;41;46m█[0m[38;2;70;69;74m█[0m[38;2;34;34;36m█[0m[38;2;70;67;62m█[0m[38;2;75;68;60m█[0m[38;2;91;78;62m█[0m[38;2;118;104;91m█[0m[38;2;147;134;118m█[0m[38;2;164;151;135m█[0m[38;2;173;161;145m█[0m[38;2;185;167;153m█[0m[38;2;193;174;160m█[0m[38;2;194;175;161m█[0m[38;2;197;178;164m█[0m[38;2;198;179;165m█[0m[38;2;200;182;168m█[0m[38;2;197;181;166m█[0m[38;2;200;184;169m█[0m[38;2;192;181;159m█[0m[38;2;183;170;151m█[0m[38;2;161;149;125m█[0m[38;2;141;131;106m█[0m[38;2;110;99;81m█[0m[38;2;73;61;47m█[0m[38;2;71;66;60m█[0m[38;2;69;61;58m█[0m[38;2;84;79;75m█[0m[38;2;71;60;58m█[0m[38;2;78;60;58m█[0m[38;2;73;56;46m█[0m[38;2;41;17;5m█[0m[38;2;73;52;33m█[0m[38;2;97;74;56m█[0m[38;2;94;73;56m█[0m[38;2;110;91;77m█[0m[38;2;100;80;69m█[0m");
$display("[38;2;0;0;0m███████████████████████████████████████[0m[38;2;1;1;1m█[0m[38;2;0;0;0m███████[0m[38;2;13;7;7m█[0m[38;2;116;98;76m█[0m[38;2;94;76;52m█[0m[38;2;76;55;34m█[0m[38;2;72;53;36m█[0m[38;2;92;70;57m█[0m[38;2;94;81;65m█[0m[38;2;106;93;77m█[0m[38;2;122;110;96m█[0m[38;2;117;109;98m█[0m[38;2;104;97;89m█[0m[38;2;60;50;49m█[0m[38;2;32;20;22m█[0m[38;2;30;22;20m█[0m[38;2;41;25;26m█[0m[38;2;51;35;36m█[0m[38;2;67;53;52m█[0m[38;2;113;98;93m█[0m[38;2;95;78;70m█[0m[38;2;103;81;68m█[0m[38;2;131;113;103m█[0m[38;2;155;136;122m█[0m[38;2;166;147;133m█[0m[38;2;175;156;142m█[0m[38;2;174;155;141m█[0m[38;2;181;162;148m█[0m[38;2;190;171;157m█[0m[38;2;193;174;160m█[0m[38;2;196;177;163m█[0m[38;2;202;180;167m█[0m[38;2;204;182;169m█[0m[38;2;204;184;173m█[0m[38;2;193;177;162m█[0m[38;2;184;160;150m█[0m[38;2;151;136;117m█[0m[38;2;106;97;80m█[0m[38;2;71;60;58m█[0m[38;2;42;41;39m█[0m[38;2;30;31;35m█[0m[38;2;22;21;26m█[0m[38;2;47;37;45m█[0m[38;2;28;21;29m█[0m[38;2;25;23;26m█[0m[38;2;30;22;19m█[0m[38;2;47;37;28m█[0m[38;2;76;64;50m█[0m[38;2;87;75;61m█[0m[38;2;76;64;48m█[0m[38;2;41;29;17m█[0m[38;2;36;26;14m█[0m");
$display("[38;2;0;0;0m█████████████████████████████████████[0m[38;2;239;235;234m█[0m[38;2;235;231;230m█[0m[38;2;206;202;201m█[0m[38;2;212;208;207m█[0m[38;2;0;0;0m█████[0m[38;2;4;0;0m█[0m[38;2;103;84;69m█[0m[38;2;107;76;55m█[0m[38;2;75;43;20m█[0m[38;2;66;40;17m█[0m[38;2;73;55;35m█[0m[38;2;96;74;60m█[0m[38;2;100;88;72m█[0m[38;2;106;94;78m█[0m[38;2;110;98;82m█[0m[38;2;131;123;102m█[0m[38;2;138;132;110m█[0m[38;2;149;143;121m█[0m[38;2;120;114;92m█[0m[38;2;99;88;68m█[0m[38;2;103;90;71m█[0m[38;2;107;92;73m█[0m[38;2;115;96;82m█[0m[38;2;110;86;74m█[0m[38;2;109;87;74m█[0m[38;2;131;112;98m█[0m[38;2;159;140;126m█[0m[38;2;167;148;134m█[0m[38;2;169;150;136m█[0m[38;2;174;155;141m██[0m[38;2;180;161;147m█[0m[38;2;191;172;158m█[0m[38;2;190;171;157m█[0m[38;2;197;178;164m██[0m[38;2;196;177;163m██[0m[38;2;190;171;157m█[0m[38;2;167;148;134m█[0m[38;2;132;113;99m█[0m[38;2;116;101;82m█[0m[38;2;78;67;63m█[0m[38;2;48;46;49m█[0m[38;2;25;25;33m█[0m[38;2;62;60;73m█[0m[38;2;92;86;96m█[0m[38;2;33;25;38m█[0m[38;2;22;20;25m█[0m[38;2;28;26;29m█[0m[38;2;43;36;26m█[0m[38;2;67;58;43m█[0m[38;2;96;89;71m█[0m[38;2;112;103;86m█[0m[38;2;108;99;82m█[0m[38;2;102;93;76m█[0m");
$display("[38;2;0;0;0m███████████████████████████████████[0m[38;2;0;1;0m█[0m[38;2;186;180;180m█[0m[38;2;213;207;207m█[0m[38;2;189;183;183m█[0m[38;2;199;190;191m█[0m[38;2;191;182;183m█[0m[38;2;90;84;86m█[0m[38;2;0;0;0m████[0m[38;2;81;66;59m█[0m[38;2;147;115;94m█[0m[38;2;110;73;47m█[0m[38;2;98;61;35m█[0m[38;2;90;55;33m█[0m[38;2;86;68;48m█[0m[38;2;113;91;77m█[0m[38;2;130;121;104m█[0m[38;2;146;137;120m█[0m[38;2;147;140;122m█[0m[38;2;154;148;126m█[0m[38;2;157;151;127m█[0m[38;2;173;167;145m█[0m[38;2;192;184;163m█[0m[38;2;204;193;173m█[0m[38;2;204;191;172m█[0m[38;2;204;189;170m█[0m[38;2;198;181;165m█[0m[38;2;188;169;155m█[0m[38;2;177;158;144m█[0m[38;2;167;148;134m█[0m[38;2;172;154;140m█[0m[38;2;173;154;140m█[0m[38;2;171;149;136m█[0m[38;2;175;151;139m█[0m[38;2;178;151;140m█[0m[38;2;189;162;151m█[0m[38;2;186;159;148m█[0m[38;2;188;161;150m█[0m[38;2;194;167;156m█[0m[38;2;199;175;163m█[0m[38;2;203;181;168m█[0m[38;2;197;178;164m█[0m[38;2;185;166;152m█[0m[38;2;145;126;112m█[0m[38;2;99;80;63m█[0m[38;2;100;81;64m█[0m[38;2;99;78;77m█[0m[38;2;104;88;89m█[0m[38;2;68;55;62m█[0m[38;2;65;47;61m█[0m[38;2;55;43;57m█[0m[38;2;37;23;38m█[0m[38;2;32;20;32m█[0m[38;2;59;47;51m█[0m[38;2;94;80;69m█[0m[38;2;106;93;77m█[0m[38;2;113;100;84m█[0m[38;2;117;106;88m█[0m[38;2;111;105;83m█[0m[38;2;96;88;65m█[0m");
$display("[38;2;0;0;0m███████████████████████████████████[0m[38;2;1;1;3m█[0m[38;2;202;195;203m█[0m[38;2;210;200;208m█[0m[38;2;195;186;189m█[0m[38;2;201;189;191m█[0m[38;2;195;186;187m█[0m[38;2;114;112;113m█[0m[38;2;0;0;0m████[0m[38;2;141;124;114m█[0m[38;2;140;110;86m█[0m[38;2;106;70;34m█[0m[38;2;89;54;22m█[0m[38;2;87;52;20m█[0m[38;2;97;71;46m█[0m[38;2;130;109;90m█[0m[38;2;146;130;115m█[0m[38;2;155;143;127m█[0m[38;2;166;159;141m█[0m[38;2;184;178;156m█[0m[38;2;198;194;169m█[0m[38;2;201;195;173m█[0m[38;2;210;203;184m█[0m[38;2;212;204;183m█[0m[38;2;209;197;175m█[0m[38;2;205;190;169m█[0m[38;2;206;189;171m█[0m[38;2;201;182;165m█[0m[38;2;200;181;164m█[0m[38;2;185;172;153m█[0m[38;2;174;155;138m█[0m[38;2;173;150;134m█[0m[38;2;167;139;125m█[0m[38;2;173;145;131m█[0m[38;2;172;144;132m█[0m[38;2;180;152;141m█[0m[38;2;187;159;148m█[0m[38;2;183;155;144m█[0m[38;2;182;154;143m█[0m[38;2;181;153;142m█[0m[38;2;191;167;155m█[0m[38;2;198;171;160m█[0m[38;2;186;168;154m█[0m[38;2;163;147;132m█[0m[38;2;147;132;113m█[0m[38;2;142;127;108m█[0m[38;2;150;134;119m█[0m[38;2;130;111;104m█[0m[38;2;106;82;78m█[0m[38;2;85;64;59m█[0m[38;2;95;71;67m█[0m[38;2;99;78;73m█[0m[38;2;116;93;85m█[0m[38;2;123;103;92m█[0m[38;2;132;113;99m█[0m[38;2;124;108;93m█[0m[38;2;123;110;94m█[0m[38;2;121;109;93m█[0m[38;2;121;113;100m█[0m[38;2;133;123;114m█[0m");
$display("[38;2;0;0;0m███████████████████████████████[0m[38;2;6;6;6m█[0m[38;2;96;96;96m█[0m[38;2;198;198;200m█[0m[38;2;212;212;214m█[0m[38;2;215;211;210m█[0m[38;2;237;231;233m█[0m[38;2;243;237;239m█[0m[38;2;224;212;212m█[0m[38;2;221;210;208m█[0m[38;2;204;200;199m█[0m[38;2;100;100;100m█[0m[38;2;0;0;0m████[0m[38;2;136;124;102m█[0m[38;2;121;97;63m█[0m[38;2;94;61;28m█[0m[38;2;79;47;9m█[0m[38;2;84;54;20m█[0m[38;2;106;84;45m█[0m[38;2;130;109;80m█[0m[38;2;145;129;106m█[0m[38;2;157;144;128m█[0m[38;2;171;159;147m█[0m[38;2;178;174;149m█[0m[38;2;180;173;155m█[0m[38;2;186;179;161m█[0m[38;2;198;189;172m█[0m[38;2;198;190;177m█[0m[38;2;196;188;167m█[0m[38;2;193;188;166m█[0m[38;2;207;188;173m█[0m[38;2;207;188;174m█[0m[38;2;204;182;168m█[0m[38;2;194;171;157m█[0m[38;2;169;146;130m█[0m[38;2;159;127;114m█[0m[38;2;160;124;112m█[0m[38;2;178;140;129m█[0m[38;2;181;147;135m█[0m[38;2;190;154;142m█[0m[38;2;198;162;148m█[0m[38;2;197;165;152m█[0m[38;2;191;159;146m█[0m[38;2;178;152;139m█[0m[38;2;186;167;153m█[0m[38;2;193;174;160m█[0m[38;2;193;171;158m█[0m[38;2;189;170;156m█[0m[38;2;199;183;168m█[0m[38;2;208;192;176m█[0m[38;2;213;197;184m█[0m[38;2;191;175;159m█[0m[38;2;182;166;150m█[0m[38;2;177;160;144m█[0m[38;2;162;140;126m█[0m[38;2;140;118;105m█[0m[38;2;130;111;94m█[0m[38;2;123;104;87m█[0m[38;2;113;98;77m█[0m[38;2;113;101;75m█[0m[38;2;115;102;85m█[0m[38;2;137;125;111m█[0m[38;2;153;143;134m█[0m[38;2;158;149;144m█[0m");
$display("[38;2;0;0;0m████████████████████████████[0m[38;2;1;1;1m█[0m[38;2;111;111;109m█[0m[38;2;227;227;227m█[0m[38;2;229;229;229m█[0m[38;2;227;227;227m█[0m[38;2;231;233;230m█[0m[38;2;227;226;221m█[0m[38;2;216;213;204m█[0m[38;2;205;202;193m█[0m[38;2;205;198;190m█[0m[38;2;177;170;162m█[0m[38;2;197;188;181m█[0m[38;2;225;224;220m█[0m[38;2;98;99;94m█[0m[38;2;0;0;2m█[0m[38;2;0;0;0m███[0m[38;2;144;128;112m█[0m[38;2;142;117;86m█[0m[38;2;140;107;76m█[0m[38;2;123;92;61m█[0m[38;2;120;89;58m█[0m[38;2;136;116;83m█[0m[38;2;145;119;92m█[0m[38;2;158;144;118m█[0m[38;2;165;149;133m█[0m[38;2;163;153;141m█[0m[38;2;168;161;143m█[0m[38;2;175;170;150m█[0m[38;2;176;169;151m█[0m[38;2;185;180;161m█[0m[38;2;188;181;162m█[0m[38;2;183;183;159m█[0m[38;2;187;181;159m█[0m[38;2;198;183;164m█[0m[38;2;206;189;173m█[0m[38;2;201;182;167m█[0m[38;2;184;162;148m█[0m[38;2;151;123;109m█[0m[38;2;148;116;103m█[0m[38;2;167;129;118m█[0m[38;2;186;139;131m█[0m[38;2;184;141;132m█[0m[38;2;192;149;140m█[0m[38;2;194;151;142m█[0m[38;2;188;154;142m█[0m[38;2;179;147;134m█[0m[38;2;170;148;134m█[0m[38;2;186;164;151m█[0m[38;2;202;183;168m█[0m[38;2;204;185;170m█[0m[38;2;211;192;178m█[0m[38;2;206;190;175m█[0m[38;2;213;200;184m█[0m[38;2;218;205;189m█[0m[38;2;211;198;182m█[0m[38;2;188;175;159m█[0m[38;2;177;161;146m█[0m[38;2;164;145;131m█[0m[38;2;140;122;108m█[0m[38;2;131;109;96m█[0m[38;2;119;104;85m█[0m[38;2;114;101;82m█[0m[38;2;114;102;78m█[0m[38;2;128;115;98m█[0m[38;2;152;142;132m█[0m[38;2;168;161;151m█[0m[38;2;180;171;166m█[0m");
$display("[38;2;0;0;0m███████████████████████████[0m[38;2;1;1;1m█[0m[38;2;236;236;236m█[0m[38;2;230;230;230m█[0m[38;2;226;226;226m█[0m[38;2;218;218;216m█[0m[38;2;209;209;197m█[0m[38;2;213;205;192m█[0m[38;2;208;205;186m█[0m[38;2;206;199;181m█[0m[38;2;194;187;169m█[0m[38;2;166;159;141m█[0m[38;2;151;139;123m█[0m[38;2;158;147;129m█[0m[38;2;183;181;166m█[0m[38;2;209;209;197m█[0m[38;2;26;27;22m█[0m[38;2;0;0;0m██[0m[38;2;2;2;4m█[0m[38;2;117;101;86m█[0m[38;2;162;132;106m█[0m[38;2;143;107;71m█[0m[38;2;124;91;56m█[0m[38;2;129;106;75m█[0m[38;2;150;133;105m█[0m[38;2;155;141;114m█[0m[38;2;168;157;135m█[0m[38;2;163;155;134m█[0m[38;2;163;156;138m█[0m[38;2;160;153;135m█[0m[38;2;161;154;136m█[0m[38;2;170;163;145m█[0m[38;2;177;172;153m█[0m[38;2;179;174;155m█[0m[38;2;174;168;152m█[0m[38;2;178;173;154m█[0m[38;2;186;178;157m█[0m[38;2;194;178;153m█[0m[38;2;193;171;148m█[0m[38;2;167;146;127m█[0m[38;2;140;108;95m█[0m[38;2;147;103;92m█[0m[38;2;166;126;118m█[0m[38;2;193;138;133m█[0m[38;2;198;148;141m█[0m[38;2;203;156;148m██[0m[38;2;176;142;130m█[0m[38;2;169;133;121m█[0m[38;2;163;137;124m█[0m[38;2;192;166;149m█[0m[38;2;216;189;172m█[0m[38;2;217;191;178m█[0m[38;2;217;196;177m█[0m[38;2;214;198;182m█[0m[38;2;213;201;185m█[0m[38;2;214;202;186m█[0m[38;2;209;197;181m█[0m[38;2;207;195;179m█[0m[38;2;201;189;173m█[0m[38;2;190;178;162m█[0m[38;2;178;162;147m█[0m[38;2;155;136;119m█[0m[38;2;142;126;110m█[0m[38;2;140;124;108m█[0m[38;2;139;132;113m█[0m[38;2;145;138;119m█[0m[38;2;160;154;132m█[0m[38;2;173;165;154m█[0m[38;2;182;173;168m█[0m");
$display("[38;2;0;0;0m██████████████████████████[0m[38;2;45;45;45m█[0m[38;2;233;233;233m█[0m[38;2;223;223;223m█[0m[38;2;223;225;222m█[0m[38;2;212;213;207m█[0m[38;2;206;208;197m█[0m[38;2;208;202;188m█[0m[38;2;204;198;176m█[0m[38;2;210;192;172m█[0m[38;2;198;181;163m█[0m[38;2;187;170;152m█[0m[38;2;158;141;123m█[0m[38;2;154;133;114m█[0m[38;2;153;132;115m█[0m[38;2;162;146;123m█[0m[38;2;182;176;152m█[0m[38;2;168;169;151m█[0m[38;2;3;3;1m█[0m[38;2;0;1;5m█[0m[38;2;1;1;3m█[0m[38;2;5;0;0m█[0m[38;2;157;135;121m█[0m[38;2;174;153;124m█[0m[38;2;172;151;124m█[0m[38;2;177;156;125m█[0m[38;2;197;175;152m█[0m[38;2;196;177;160m█[0m[38;2;192;179;163m█[0m[38;2;184;171;155m█[0m[38;2;177;165;149m█[0m[38;2;170;161;144m█[0m[38;2;158;151;133m█[0m[38;2;159;152;134m█[0m[38;2;166;159;141m█[0m[38;2;171;164;146m█[0m[38;2;174;167;149m█[0m[38;2;172;164;143m█[0m[38;2;176;166;141m█[0m[38;2;183;167;142m█[0m[38;2;183;161;138m█[0m[38;2;163;143;119m█[0m[38;2;154;119;100m█[0m[38;2;167;119;105m█[0m[38;2;151;109;93m█[0m[38;2;168;114;102m█[0m[38;2;178;129;115m█[0m[38;2;180;134;119m█[0m[38;2;179;133;118m█[0m[38;2;170;128;112m█[0m[38;2;173;134;117m█[0m[38;2;172;141;121m█[0m[38;2;186;159;138m█[0m[38;2;211;185;162m█[0m[38;2;205;183;159m█[0m[38;2;200;179;160m█[0m[38;2;196;178;164m█[0m[38;2;194;185;168m█[0m[38;2;193;184;167m█[0m[38;2;192;183;166m█[0m[38;2;198;189;172m█[0m[38;2;197;188;171m█[0m[38;2;190;181;164m█[0m[38;2;180;171;154m█[0m[38;2;157;148;131m█[0m[38;2;152;143;126m█[0m[38;2;158;149;132m█[0m[38;2;154;147;129m█[0m[38;2;164;157;139m█[0m[38;2;169;163;139m█[0m[38;2;177;171;149m█[0m[38;2;187;177;175m█[0m");
$display("[38;2;0;0;0m████████████████████████[0m[38;2;1;1;1m█[0m[38;2;21;21;21m█[0m[38;2;242;238;239m█[0m[38;2;233;229;230m█[0m[38;2;204;200;199m█[0m[38;2;189;185;184m█[0m[38;2;175;172;165m█[0m[38;2;167;158;149m█[0m[38;2;176;161;142m█[0m[38;2;177;161;136m█[0m[38;2;182;154;132m█[0m[38;2;177;146;118m█[0m[38;2;172;142;114m█[0m[38;2;167;136;108m█[0m[38;2;154;120;93m█[0m[38;2;156;122;95m█[0m[38;2;166;136;112m█[0m[38;2;179;152;131m█[0m[38;2;185;162;146m█[0m[38;2;6;2;1m█[0m[38;2;1;0;5m█[0m[38;2;1;0;0m█[0m[38;2;1;1;3m█[0m[38;2;122;105;95m█[0m[38;2;194;177;151m█[0m[38;2;191;173;149m█[0m[38;2;198;181;155m█[0m[38;2;201;181;157m█[0m[38;2;197;179;159m█[0m[38;2;199;183;167m█[0m[38;2;190;177;160m█[0m[38;2;187;171;156m█[0m[38;2;168;156;140m█[0m[38;2;164;155;138m█[0m[38;2;155;143;127m█[0m[38;2;158;149;132m█[0m[38;2;157;148;131m█[0m[38;2;163;154;137m█[0m[38;2;169;161;142m█[0m[38;2;175;164;144m█[0m[38;2;182;167;146m█[0m[38;2;185;162;144m█[0m[38;2;170;144;127m█[0m[38;2;172;139;124m█[0m[38;2;181;133;123m█[0m[38;2;147;105;93m█[0m[38;2;150;100;91m█[0m[38;2;143;95;85m█[0m[38;2;159;112;102m█[0m[38;2;174;127;117m█[0m[38;2;192;150;136m█[0m[38;2;187;147;135m█[0m[38;2;186;153;138m█[0m[38;2;187;160;141m█[0m[38;2;196;169;150m█[0m[38;2;195;173;152m█[0m[38;2;193;172;155m█[0m[38;2;189;171;157m█[0m[38;2;187;174;158m██[0m[38;2;190;177;161m█[0m[38;2;191;179;163m█[0m[38;2;189;180;163m█[0m[38;2;181;174;156m█[0m[38;2;170;161;144m█[0m[38;2;169;160;143m█[0m[38;2;167;158;141m█[0m[38;2;169;160;143m█[0m[38;2;172;165;147m█[0m[38;2;177;170;152m█[0m[38;2;179;173;151m█[0m[38;2;181;174;155m█[0m[38;2;179;170;161m█[0m");
$display("[38;2;0;0;0m█████████████████████████[0m[38;2;170;169;167m█[0m[38;2;213;209;208m█[0m[38;2;213;203;204m█[0m[38;2;205;195;196m█[0m[38;2;208;198;197m█[0m[38;2;201;193;182m█[0m[38;2;198;193;173m█[0m[38;2;203;190;171m█[0m[38;2;189;175;149m█[0m[38;2;171;146;124m█[0m[38;2;167;136;108m█[0m[38;2;159;128;100m█[0m[38;2;149;118;90m█[0m[38;2;146;114;89m█[0m[38;2;162;130;105m█[0m[38;2;167;135;110m█[0m[38;2;169;142;121m█[0m[38;2;175;153;139m█[0m[38;2;70;64;52m█[0m[38;2;0;0;2m█[0m[38;2;2;0;1m█[0m[38;2;0;1;3m█[0m[38;2;124;111;102m█[0m[38;2;196;179;153m█[0m[38;2;204;187;159m█[0m[38;2;202;185;157m█[0m[38;2;202;185;159m█[0m[38;2;201;183;161m█[0m[38;2;198;179;162m█[0m[38;2;198;175;159m█[0m[38;2;187;169;155m█[0m[38;2;180;167;151m█[0m[38;2;168;155;139m█[0m[38;2;162;146;131m█[0m[38;2;164;148;133m█[0m[38;2;165;149;134m█[0m[38;2;163;147;132m█[0m[38;2;159;143;128m█[0m[38;2;163;150;134m█[0m[38;2;156;149;133m█[0m[38;2;163;140;132m█[0m[38;2;156;129;120m█[0m[38;2;158;123;117m█[0m[38;2;162;114;114m█[0m[38;2;159;113;113m█[0m[38;2;159;109;110m█[0m[38;2;153;103;104m█[0m[38;2;166;118;118m█[0m[38;2;167;119;119m█[0m[38;2;176;136;134m█[0m[38;2;179;141;138m█[0m[38;2;178;149;143m█[0m[38;2;186;157;151m█[0m[38;2;190;161;155m█[0m[38;2;185;161;149m█[0m[38;2;185;163;150m█[0m[38;2;187;169;155m█[0m[38;2;185;172;156m█[0m[38;2;184;171;155m█[0m[38;2;186;173;157m█[0m[38;2;188;175;159m█[0m[38;2;188;176;160m█[0m[38;2;180;173;155m█[0m[38;2;167;160;142m█[0m[38;2;171;164;146m█[0m[38;2;178;171;153m█[0m[38;2;180;173;155m█[0m[38;2;179;172;154m█[0m[38;2;179;172;156m█[0m[38;2;176;169;151m█[0m[38;2;177;170;154m█[0m[38;2;178;169;162m█[0m");
$display("[38;2;0;0;0m█████████████████████████[0m[38;2;153;159;155m█[0m[38;2;211;213;210m█[0m[38;2;208;205;200m█[0m[38;2;204;190;187m█[0m[38;2;204;186;182m█[0m[38;2;203;186;179m█[0m[38;2;196;179;171m█[0m[38;2;194;177;167m█[0m[38;2;196;173;159m█[0m[38;2;188;162;149m█[0m[38;2;172;144;123m█[0m[38;2;152;124;100m█[0m[38;2;147;119;97m█[0m[38;2;158;130;108m█[0m[38;2;162;134;113m█[0m[38;2;164;140;114m█[0m[38;2;161;140;113m█[0m[38;2;165;151;125m█[0m[38;2;153;147;131m█[0m[38;2;42;43;38m█[0m[38;2;2;0;3m█[0m[38;2;2;2;2m█[0m[38;2;123;114;109m█[0m[38;2;206;189;171m█[0m[38;2;202;190;166m█[0m[38;2;206;190;165m█[0m[38;2;208;191;163m█[0m[38;2;205;188;160m█[0m[38;2;203;186;160m█[0m[38;2;199;181;159m█[0m[38;2;194;178;152m█[0m[38;2;185;169;154m█[0m[38;2;184;171;155m█[0m[38;2;171;158;142m█[0m[38;2;168;155;139m█[0m[38;2;164;146;132m█[0m[38;2;163;141;128m██[0m[38;2;163;142;125m█[0m[38;2;161;143;123m█[0m[38;2;153;135;115m█[0m[38;2;146;133;114m█[0m[38;2;147;120;109m█[0m[38;2;149;119;109m█[0m[38;2;149;115;106m█[0m[38;2;152;113;106m█[0m[38;2;150;107;101m█[0m[38;2;152;113;106m█[0m[38;2;139;109;99m█[0m[38;2;146;119;108m█[0m[38;2;160;132;121m█[0m[38;2;169;141;130m█[0m[38;2;176;148;137m█[0m[38;2;178;150;139m█[0m[38;2;174;150;138m█[0m[38;2;177;153;141m█[0m[38;2;179;160;146m█[0m[38;2;182;160;147m█[0m[38;2;185;163;150m█[0m[38;2;186;167;153m█[0m[38;2;176;160;145m█[0m[38;2;165;152;136m█[0m[38;2;156;151;132m█[0m[38;2;164;157;138m█[0m[38;2;163;157;133m█[0m[38;2;162;156;134m█[0m[38;2;162;154;141m█[0m[38;2;157;148;139m█[0m[38;2;156;147;140m█[0m[38;2;160;151;144m█[0m[38;2;174;165;158m█[0m[38;2;170;160;158m█[0m");
$display("[38;2;0;0;0m█████████████████████████[0m[38;2;11;11;13m█[0m[38;2;232;227;223m█[0m[38;2;198;189;184m█[0m[38;2;184;169;162m█[0m[38;2;183;169;160m█[0m[38;2;177;169;150m█[0m[38;2;179;161;147m█[0m[38;2;172;153;136m█[0m[38;2;171;148;132m█[0m[38;2;176;148;134m█[0m[38;2;165;135;111m█[0m[38;2;155;124;103m█[0m[38;2;160;129;108m█[0m[38;2;154;126;104m█[0m[38;2;155;127;106m█[0m[38;2;149;125;99m█[0m[38;2;150;133;105m█[0m[38;2;161;147;118m█[0m[38;2;175;165;140m█[0m[38;2;186;181;162m█[0m[38;2;196;194;179m█[0m[38;2;145;136;127m█[0m[38;2;95;87;76m█[0m[38;2;163;155;136m█[0m[38;2;192;180;156m█[0m[38;2;198;185;166m█[0m[38;2;204;186;166m█[0m[38;2;201;183;163m█[0m[38;2;196;178;156m█[0m[38;2;195;176;159m█[0m[38;2;206;185;166m█[0m[38;2;202;188;177m█[0m[38;2;205;187;173m█[0m[38;2;195;179;164m█[0m[38;2;193;177;162m█[0m[38;2;178;156;143m█[0m[38;2;166;150;134m█[0m[38;2;164;143;122m█[0m[38;2;160;136;112m█[0m[38;2;160;134;111m█[0m[38;2;161;133;111m█[0m[38;2;157;133;121m█[0m[38;2;149;123;110m█[0m[38;2;150;123;112m█[0m[38;2;153;134;120m█[0m[38;2;155;128;117m█[0m[38;2;155;131;119m█[0m[38;2;152;128;116m█[0m[38;2;146;124;111m█[0m[38;2;146;119;108m█[0m[38;2;153;125;114m█[0m[38;2;161;133;122m█[0m[38;2;166;138;127m█[0m[38;2;172;144;133m█[0m[38;2;167;143;131m█[0m[38;2;168;146;133m█[0m[38;2;171;149;136m█[0m[38;2;169;150;136m█[0m[38;2;168;149;135m█[0m[38;2;159;143;128m█[0m[38;2;149;140;123m█[0m[38;2;146;139;121m█[0m[38;2;151;144;126m█[0m[38;2;164;157;139m█[0m[38;2;169;162;144m█[0m[38;2;181;174;156m█[0m[38;2;180;172;161m█[0m[38;2;179;170;161m█[0m[38;2;178;169;160m██[0m[38;2;179;170;161m█[0m[38;2;184;175;170m█[0m");
$display("[38;2;0;0;0m█████████████████████████[0m[38;2;0;0;2m█[0m[38;2;118;110;107m█[0m[38;2;198;188;179m█[0m[38;2;182;170;154m█[0m[38;2;179;163;140m█[0m[38;2;175;164;134m█[0m[38;2;168;156;130m█[0m[38;2;167;147;120m█[0m[38;2;157;133;109m█[0m[38;2;166;135;114m█[0m[38;2;165;133;112m█[0m[38;2;159;128;107m█[0m[38;2;162;131;110m█[0m[38;2;160;132;110m█[0m[38;2;159;131;109m█[0m[38;2;155;123;102m█[0m[38;2;164;138;113m█[0m[38;2;173;149;123m█[0m[38;2;175;159;126m█[0m[38;2;180;165;144m█[0m[38;2;179;170;155m█[0m[38;2;204;194;185m█[0m[38;2;225;215;205m█[0m[38;2;211;203;184m█[0m[38;2;179;168;150m█[0m[38;2;189;176;160m█[0m[38;2;202;183;169m█[0m[38;2;212;190;177m█[0m[38;2;208;186;175m█[0m[38;2;204;184;173m█[0m[38;2;206;187;173m██[0m[38;2;204;185;171m█[0m[38;2;198;179;165m█[0m[38;2;199;180;165m█[0m[38;2;194;176;162m█[0m[38;2;180;165;144m█[0m[38;2;168;152;127m█[0m[38;2;166;141;119m█[0m[38;2;171;145;118m█[0m[38;2;169;143;120m█[0m[38;2;184;156;144m█[0m[38;2;189;159;151m█[0m[38;2;184;155;151m█[0m[38;2;180;152;148m█[0m[38;2;175;145;134m█[0m[38;2;169;150;135m█[0m[38;2;169;145;133m█[0m[38;2;164;140;128m█[0m[38;2;162;135;124m██[0m[38;2;162;134;123m█[0m[38;2;162;132;122m█[0m[38;2;159;131;120m█[0m[38;2;159;135;123m█[0m[38;2;164;142;129m█[0m[38;2;162;140;127m█[0m[38;2;152;133;119m█[0m[38;2;155;136;122m█[0m[38;2;156;140;125m█[0m[38;2;166;153;137m█[0m[38;2;167;155;141m█[0m[38;2;164;158;142m█[0m[38;2;167;161;139m█[0m[38;2;178;171;153m█[0m[38;2;180;173;157m█[0m[38;2;176;168;155m█[0m[38;2;178;169;160m█[0m[38;2;176;167;158m█[0m[38;2;188;179;170m█[0m[38;2;189;180;171m█[0m[38;2;189;179;177m█[0m");
$display("[38;2;0;0;0m██████████████████████████[0m[38;2;1;1;1m█[0m[38;2;66;65;61m█[0m[38;2;170;165;159m█[0m[38;2;188;181;171m█[0m[38;2;177;170;154m█[0m[38;2;176;163;147m█[0m[38;2;169;153;130m█[0m[38;2;163;147;122m█[0m[38;2;170;143;122m█[0m[38;2;170;148;124m█[0m[38;2;160;138;114m█[0m[38;2;162;140;116m█[0m[38;2;162;136;113m█[0m[38;2;166;140;117m█[0m[38;2;168;142;119m█[0m[38;2;177;149;127m█[0m[38;2;185;159;136m█[0m[38;2;179;159;134m█[0m[38;2;181;160;139m█[0m[38;2;184;167;147m█[0m[38;2;191;178;162m█[0m[38;2;202;189;173m█[0m[38;2;201;188;172m█[0m[38;2;206;193;177m█[0m[38;2;193;180;164m█[0m[38;2;197;184;168m█[0m[38;2;204;191;175m█[0m[38;2;203;190;174m█[0m[38;2;204;191;175m█[0m[38;2;205;186;172m█[0m[38;2;206;187;173m█[0m[38;2;202;183;169m█[0m[38;2;199;180;166m█[0m[38;2;198;179;164m█[0m[38;2;197;179;165m█[0m[38;2;193;179;153m█[0m[38;2;189;169;145m█[0m[38;2;186;162;138m█[0m[38;2;183;157;134m█[0m[38;2;186;160;137m█[0m[38;2;183;159;135m██[0m[38;2;181;155;132m█[0m[38;2;180;152;130m█[0m[38;2;184;157;138m█[0m[38;2;183;157;144m█[0m[38;2;185;158;147m█[0m[38;2;181;154;143m█[0m[38;2;184;156;145m█[0m[38;2;186;158;147m██[0m[38;2;187;159;148m█[0m[38;2;182;154;143m█[0m[38;2;172;148;136m█[0m[38;2;172;150;137m█[0m[38;2;175;153;140m█[0m[38;2;175;156;142m█[0m[38;2;174;155;141m█[0m[38;2;167;149;137m█[0m[38;2;169;153;140m█[0m[38;2;173;159;148m█[0m[38;2;174;165;156m█[0m[38;2;175;166;157m█[0m[38;2;176;167;158m█[0m[38;2;178;169;160m█[0m[38;2;181;172;163m█[0m[38;2;180;171;162m█[0m[38;2;182;173;164m█[0m[38;2;177;168;159m██[0m[38;2;180;170;168m█[0m");
$display("[38;2;0;0;0m█████████████████████████████[0m[38;2;1;3;2m█[0m[38;2;139;131;129m█[0m[38;2;191;180;176m█[0m[38;2;189;175;166m█[0m[38;2;188;172;156m█[0m[38;2;182;161;140m█[0m[38;2;168;152;126m█[0m[38;2;170;153;127m█[0m[38;2;173;151;127m█[0m[38;2;174;150;126m█[0m[38;2;181;155;132m█[0m[38;2;185;159;136m█[0m[38;2;191;163;141m█[0m[38;2;185;161;137m█[0m[38;2;185;163;139m█[0m[38;2;180;158;134m█[0m[38;2;189;168;141m█[0m[38;2;183;166;138m█[0m[38;2;195;176;159m█[0m[38;2;189;170;156m█[0m[38;2;199;180;166m█[0m[38;2;212;190;177m█[0m[38;2;196;183;167m█[0m[38;2;190;177;161m█[0m[38;2;192;179;163m█[0m[38;2;201;188;172m█[0m[38;2;203;184;170m█[0m[38;2;205;186;172m█[0m[38;2;201;182;168m█[0m[38;2;202;183;169m██[0m[38;2;198;179;165m█[0m[38;2;196;180;154m█[0m[38;2;187;167;142m█[0m[38;2;186;162;138m█[0m[38;2;181;157;133m█[0m[38;2;177;153;129m█[0m[38;2;176;151;120m█[0m[38;2;175;149;122m█[0m[38;2;172;146;119m█[0m[38;2;174;148;121m█[0m[38;2;171;146;116m█[0m[38;2;165;139;114m█[0m[38;2;174;148;123m█[0m[38;2;182;156;131m█[0m[38;2;185;158;139m█[0m[38;2;177;150;131m██[0m[38;2;173;147;132m█[0m[38;2;177;152;132m█[0m[38;2;171;146;126m█[0m[38;2;175;148;131m█[0m[38;2;168;151;135m█[0m[38;2;169;150;135m█[0m[38;2;167;147;136m█[0m[38;2;164;148;133m█[0m[38;2;173;159;146m█[0m[38;2;169;159;147m█[0m[38;2;169;159;150m█[0m[38;2;165;155;146m█[0m[38;2;164;157;147m█[0m[38;2;165;156;147m█[0m[38;2;163;154;145m█[0m[38;2;161;157;146m█[0m[38;2;165;163;151m█[0m[38;2;169;167;155m█[0m[38;2;176;172;161m█[0m[38;2;174;166;163m█[0m");
$display("[38;2;0;0;0m███████████████████████████████[0m[38;2;217;216;212m█[0m[38;2;209;202;194m█[0m[38;2;203;195;182m█[0m[38;2;199;186;169m█[0m[38;2;178;171;143m█[0m[38;2;177;163;137m█[0m[38;2;178;160;136m█[0m[38;2;189;165;139m█[0m[38;2;186;158;136m█[0m[38;2;193;167;144m█[0m[38;2;191;167;143m█[0m[38;2;186;162;138m█[0m[38;2;188;162;139m█[0m[38;2;193;167;144m█[0m[38;2;185;163;140m█[0m[38;2;189;171;147m█[0m[38;2;187;168;151m█[0m[38;2;183;164;150m█[0m[38;2;194;175;161m█[0m[38;2;195;179;164m█[0m[38;2;199;186;170m█[0m[38;2;188;175;159m█[0m[38;2;183;170;154m█[0m[38;2;175;162;146m█[0m[38;2;193;177;162m█[0m[38;2;204;182;169m█[0m[38;2;191;173;159m█[0m[38;2;193;174;160m█[0m[38;2;195;176;162m█[0m[38;2;194;175;161m█[0m[38;2;195;178;152m█[0m[38;2;194;177;151m█[0m[38;2;194;174;149m█[0m[38;2;194;170;146m█[0m[38;2;183;159;135m█[0m[38;2;178;152;125m█[0m[38;2;174;148;113m█[0m[38;2;169;144;113m█[0m[38;2;167;142;111m█[0m[38;2;162;137;107m█[0m[38;2;169;144;114m█[0m[38;2;174;149;119m█[0m[38;2;176;151;121m█[0m[38;2;169;144;114m█[0m[38;2;165;140;110m█[0m[38;2;171;148;117m█[0m[38;2;164;140;114m█[0m[38;2;168;144;118m█[0m[38;2;175;151;125m█[0m[38;2;169;148;119m█[0m[38;2;163;140;122m█[0m[38;2;164;146;126m█[0m[38;2;169;150;135m█[0m[38;2;164;145;130m█[0m[38;2;162;145;137m█[0m[38;2;154;144;134m█[0m[38;2;153;138;133m█[0m[38;2;145;135;126m█[0m[38;2;136;126;117m█[0m[38;2;135;126;117m█[0m[38;2;136;127;118m█[0m[38;2;128;126;114m█[0m[38;2;134;130;119m█[0m[38;2;137;133;122m█[0m[38;2;143;139;128m█[0m[38;2;145;140;134m█[0m");
$display("[38;2;0;0;0m███████████████████████████████[0m[38;2;2;2;2m█[0m[38;2;224;224;226m█[0m[38;2;213;218;214m█[0m[38;2;206;203;194m█[0m[38;2;189;182;166m█[0m[38;2;182;170;156m█[0m[38;2;178;161;151m█[0m[38;2;186;164;143m█[0m[38;2;185;162;144m█[0m[38;2;193;166;145m█[0m[38;2;193;167;144m██[0m[38;2;186;158;136m█[0m[38;2;189;161;139m█[0m[38;2;188;166;143m█[0m[38;2;187;168;153m█[0m[38;2;184;165;148m█[0m[38;2;180;161;147m█[0m[38;2;192;170;157m█[0m[38;2;188;170;156m█[0m[38;2;189;176;160m██[0m[38;2;187;178;161m█[0m[38;2;188;185;166m█[0m[38;2;191;175;160m█[0m[38;2;190;171;157m█[0m[38;2;196;177;163m█[0m[38;2;197;178;163m█[0m[38;2;199;179;168m█[0m[38;2;198;179;162m█[0m[38;2;193;175;151m██[0m[38;2;196;176;151m█[0m[38;2;194;170;146m█[0m[38;2;186;162;138m█[0m[38;2;181;156;126m█[0m[38;2;176;150;117m█[0m[38;2;174;150;114m█[0m[38;2;160;136;98m█[0m[38;2;163;138;108m█[0m[38;2;166;141;111m█[0m[38;2;167;142;112m█[0m[38;2;166;141;111m█[0m[38;2;176;151;120m█[0m[38;2;182;156;129m█[0m[38;2;178;154;128m█[0m[38;2;182;157;135m█[0m[38;2;174;150;126m█[0m[38;2;168;142;119m█[0m[38;2;169;143;120m█[0m[38;2;156;135;106m█[0m[38;2;153;136;110m█[0m[38;2;139;120;103m█[0m[38;2;139;121;101m█[0m[38;2;140;124;111m█[0m[38;2;135;117;113m█[0m[38;2;141;124;116m█[0m[38;2;143;123;114m█[0m[38;2;122;109;101m█[0m[38;2;113;104;95m█[0m[38;2;108;99;90m█[0m[38;2;101;97;86m█[0m[38;2;105;101;92m█[0m[38;2;121;117;106m█[0m[38;2;126;122;111m█[0m[38;2;130;125;121m█[0m");
$display("[38;2;0;0;0m████████████████████████████████[0m[38;2;48;48;48m█[0m[38;2;211;213;212m█[0m[38;2;204;206;205m█[0m[38;2;191;197;183m█[0m[38;2;189;185;173m█[0m[38;2;185;179;157m█[0m[38;2;191;177;148m█[0m[38;2;192;170;146m█[0m[38;2;196;172;148m█[0m[38;2;189;171;147m█[0m[38;2;189;172;146m█[0m[38;2;187;169;149m█[0m[38;2;188;170;150m█[0m[38;2;188;169;155m█[0m[38;2;187;168;154m█[0m[38;2;185;166;152m█[0m[38;2;173;154;140m█[0m[38;2;186;164;151m█[0m[38;2;185;167;153m█[0m[38;2;184;171;155m█[0m[38;2;188;175;159m██[0m[38;2;187;174;158m█[0m[38;2;183;167;154m█[0m[38;2;179;159;148m█[0m[38;2;194;175;161m█[0m[38;2;198;181;163m█[0m[38;2;197;181;165m█[0m[38;2;195;178;162m█[0m[38;2;196;177;162m█[0m[38;2;192;173;158m█[0m[38;2;195;174;157m█[0m[38;2;196;170;153m█[0m[38;2;197;171;154m█[0m[38;2;191;164;145m█[0m[38;2;191;163;142m█[0m[38;2;183;157;134m█[0m[38;2;186;160;135m█[0m[38;2;184;158;135m█[0m[38;2;168;145;113m█[0m[38;2;169;146;115m█[0m[38;2;166;143;112m█[0m[38;2;165;139;112m█[0m[38;2;166;140;113m█[0m[38;2;161;137;113m█[0m[38;2;168;144;118m█[0m[38;2;162;136;113m█[0m[38;2;152;130;106m█[0m[38;2;141;121;96m█[0m[38;2;137;120;90m█[0m[38;2;125;111;82m█[0m[38;2;121;106;85m█[0m[38;2;121;100;79m█[0m[38;2;118;96;85m█[0m[38;2;109;91;89m█[0m[38;2;124;106;104m█[0m[38;2;118;103;100m█[0m[38;2;93;82;78m█[0m[38;2;91;82;73m█[0m[38;2;81;72;63m█[0m[38;2;82;78;69m█[0m[38;2;80;75;69m█[0m[38;2;87;82;76m█[0m[38;2;94;89;83m█[0m[38;2;96;91;85m█[0m");
$display("[38;2;0;0;0m████████████████████████████████[0m[38;2;19;19;19m█[0m[38;2;206;206;206m█[0m[38;2;194;194;194m█[0m[38;2;191;193;180m█[0m[38;2;192;182;170m█[0m[38;2;194;179;160m█[0m[38;2;187;169;145m█[0m[38;2;200;169;149m█[0m[38;2;196;169;148m█[0m[38;2;195;173;150m█[0m[38;2;196;174;151m█[0m[38;2;190;165;145m█[0m[38;2;194;169;149m█[0m[38;2;191;170;153m█[0m[38;2;188;169;155m█[0m[38;2;185;166;151m█[0m[38;2;182;163;148m█[0m[38;2;182;160;146m█[0m[38;2;183;166;150m██[0m[38;2;181;164;148m██[0m[38;2;183;166;150m█[0m[38;2;181;164;146m█[0m[38;2;189;166;148m█[0m[38;2;194;171;153m█[0m[38;2;194;172;149m█[0m[38;2;192;172;148m█[0m[38;2;190;168;147m█[0m[38;2;190;165;145m█[0m[38;2;185;163;142m█[0m[38;2;193;168;148m█[0m[38;2;192;165;146m█[0m[38;2;189;164;144m█[0m[38;2;191;164;143m█[0m[38;2;189;163;140m█[0m[38;2;188;162;137m█[0m[38;2;184;158;135m█[0m[38;2;187;160;139m█[0m[38;2;179;155;129m█[0m[38;2;180;156;128m█[0m[38;2;175;151;123m█[0m[38;2;175;149;124m█[0m[38;2;172;148;122m█[0m[38;2;168;146;122m█[0m[38;2;168;147;120m█[0m[38;2;164;144;119m█[0m[38;2;160;144;118m█[0m[38;2;142;128;102m█[0m[38;2;132;121;101m█[0m[38;2;112;101;83m█[0m[38;2;109;99;87m█[0m[38;2;103;91;75m█[0m[38;2;87;77;67m█[0m[38;2;84;73;69m█[0m[38;2;80;69;67m█[0m[38;2;70;56;53m█[0m[38;2;48;37;35m█[0m[38;2;49;39;37m██[0m[38;2;46;39;33m█[0m[38;2;51;44;38m█[0m[38;2;63;56;50m█[0m[38;2;62;55;49m█[0m[38;2;54;49;43m█[0m");
$display("\n");
$display("                              \033[32m\033[5m █████ █████ █████ █████ █████ █████ █████ \033[0m");
$display("                              \033[32m\033[5m █     █   █ █   █ █   █ █     █       █ \033[0m");
$display("                              \033[32m\033[5m █     █   █ █████ █████ █████ █       █  \033[0m");
$display("                              \033[32m\033[5m █     █   █ █  █  █  █  █     █       █  \033[0m");
$display("                              \033[32m\033[5m █████ █████ █   █ █   █ █████ █████   █  \033[0m");
$display("\n");

end endtask

endmodule
