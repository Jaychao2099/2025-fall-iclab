`ifdef FUNC
`define LAT_MAX 20
`define LAT_MIN 1
`endif
`ifdef PERF
`define LAT_MAX 500
`define LAT_MIN 300
`endif

module pseudo_DRAM_data#(parameter ID_WIDTH=4, ADDR_WIDTH=32, DATA_WIDTH=16, BURST_LEN=7) (
// Glbal Signal
  	  input clk,
  	  input rst_n,
// slave interface 
      // axi write address channel 
      // src master
      input wire [ID_WIDTH-1:0]     awid_s_inf,
      input wire [ADDR_WIDTH-1:0] awaddr_s_inf,
      input wire [2:0]            awsize_s_inf,
      input wire [1:0]           awburst_s_inf,
      input wire [BURST_LEN-1:0]   awlen_s_inf,
      input wire                 awvalid_s_inf,
      // src slave
      output reg                 awready_s_inf,
      // -----------------------------
   
      // axi write data channel 
      // src master
      input wire [DATA_WIDTH-1:0]  wdata_s_inf,
      input wire                   wlast_s_inf,
      input wire                  wvalid_s_inf,
      // src slave
      output reg                  wready_s_inf,
   
      // axi write response channel 
      // src slave
      output reg  [ID_WIDTH-1:0]     bid_s_inf,
      output reg  [1:0]            bresp_s_inf,
      output reg                  bvalid_s_inf,
      // src master 
      input wire                  bready_s_inf,
      // -----------------------------
   
      // axi read address channel 
      // src master
      input wire [ID_WIDTH-1:0]     arid_s_inf,
      input wire [ADDR_WIDTH-1:0] araddr_s_inf,
      input wire [BURST_LEN-1:0]   arlen_s_inf,
      input wire [2:0]            arsize_s_inf,
      input wire [1:0]           arburst_s_inf,
      input wire                 arvalid_s_inf,
      // src slave
      output reg                 arready_s_inf,
      // -----------------------------
   
      // axi read data channel 
      // slave
      output reg [ID_WIDTH-1:0]      rid_s_inf,
      output reg [DATA_WIDTH-1:0]  rdata_s_inf,
      output reg [1:0]             rresp_s_inf,
      output reg                   rlast_s_inf,
      output reg                  rvalid_s_inf,
      // master
      input wire                  rready_s_inf
      // -----------------------------
);

`protected
NNKWQ6FBg5)Pf&WG<]2;P:,]5gQSDNIWf&DM=_<:@d6e7#6f+1M/0)S+17H4IIZ7
RD54#=UIZQ>MT&OaMYe^7-ZG#YK5dVFHfQ].6Y#NP/#GfF.:aDXV7PRC&B#a\]1[
dU5d3[\PUYS(&O,N[X@\gf3ZV9IN0)b;=Z0;GR=V.1:1@BCZG@:..AL^.S8H>9OM
B)/c&<eW&\,[aR8;H8<;FO=0f4VTBXW-M6#,7Jb^CS<G?OHWF2WFbTeQ11^gD)[_
6G(/>ceb0FI41f&(7(9P&N<^9BMTT>?P0,E_TaDBGg8O/=H:SI?A(T@8]aSRD)BW
FNeDaFI\S[ZB&<F<=6P)AT,B-9#UBFKJg(<-RQ^7acWaAJNM1O^Ia?g?:))Y[OL/
Y,GXL<FDe]\Z._9,5E+J4UU7R>bMEDVY[Q^/23OW(P+\Tb\X:KH=E7UV-D_cP)9B
LNb23dEXAI7;].,McSMHN((;&3+J&8O0O,[J+c0@O\F2aBV/4A#CbbGR3K&8OKX<
=H\bNK1C?_b13<9GDEARR9_,L7VWAX51P-R[5^]>@X>]B:H5H[8LJ;,D2ELJRaA[
+P.<+#MCb)D?a[T+#PVa[F1BPZ+7D-<T)-)b1X07MREg?_0d.HQ<FNYL&;5MdFQ@
:^.\D4#KDVff+\#XZGRTAFHC.A[(I60D6Fa>dDKOZQeI?bXDJ4eLQb?U]11Q@X80
@\#_g_X1+Pe23@f.6A8=L(QCY@Of,/(4Z=D-9BFdI/S^59fEF\/B432gDfOLD6DC
Se1Y)(5R940eJMRE7H,I+/]:f&@8Q<]M[[/W5O9N(,HD,@+f-c_eA0:E9/Y0gOD-
Be7CQEHYBOYFgP_)1D&B([U^B:+Wd4^6_a@?CUQ8M2#F])K9_Z4B1;Hg[B#LZ6U#
_799\M0(\L,:/=Pd.>LDB8:f,KM6H@UX39GTCHb4&6QD/.,[Q.@Nf5WXUFe8d(f-
:;1NH_cfEUd,E[B3.c1S,A^dFNI\6]Gc5@+;6f19SP3f^5;?WTc8Q\JG14&X8Q7K
&2]4BG9+T2ZMFD(KEB8cH2dHQ]QTMCN\H+SU&8e][W?8Sa?:7@0T-?0Q,5;,Y4GY
9Ma)UM>A@_P;Q)<6a+C8U><ZfJT#bKM)0-=_[#aRJ;J\=BAc:J=FEKMQ7K<E:&VD
&GDFGdXDaI2K0^.[6_9&=KZ\CM3-L;>2+<14-\fKEN\:G8UY_)\H3Z?<]@gT1S.e
a(UA&/fGH,&LQe04f-Ne)KB=M??ABX3Z6f42WE#5.&(M@XQ.&K2O:NS+g<4??)ZB
d#5C.##K,D76;:YgYQPQ<K\;:7R9.Y;8dB9W1KX4L[1&U?)g;H;PYBAEH6[4<L\/
]Q2a\G>GFX-<]4>066?4N2Z)Q7:#B;NSR+?f=?42dS4C1VG2<)L+G68:I3J8a<XL
F@?N7/W<>NC58>AgT\IB.e48<LR5f>IC7b=.8/2/-E&7(=O>8(+T(PD<fbKAWP=O
gb4(_.VN<^F2N#&IbZ.S6W+;ca(LSM+-O5A9/c=UC_TeA&B&b-N-e4(,BWe<]EBB
G5&(X_W&,@#XR#K6GR8MQPd>=S9W^;UXcfRJcL^0;<MW-NHbW^W86YY>G[1UZZAM
4,JUFee#J\.Rb1;-2\^:fT0L+64e_&@NA9Va;P6DT.?PR,VGIgGf&MX5J<W4d6Z&
aR8J-2:M/PH+U-2,J)P0\Z2QeP362bR#FZNN38N^])166:?/)B4>MVRW.-GBIRBg
(N#02CGP^BDVb^P>C21#1978UJ4AN4DVLRHAfOC9=HI\UY-dC[(^6&\O4geH(6[.
WG^R@-S71Rb0c.5B76(c:DA)Q3:E@;;N>3NDPaK.&VW;O.E<#W6OEH>(5DbDM-Lb
[,#cCQaS&8e=MAFU.?UcIgT1[20QDSH_50X][DcgY#L/:&N>c)?c<+3@PPgSEFBB
UECVLbO_[d71(9UK_,F?cAKW;XL>22NMcTQ.8gdSLI8&(D1--[/B55ZHc=4D6SAV
3?U)HP1V))_@K6gF-][\;[=&OcfYDIF9e4NEUA&d4N#47ZSEYY6fMI=-Z/:X2G,f
9YDP<JfgR5-,OY8+RT4UPZ;##f:&b=MMQFD03A>PbgW/R57gTd=-aV-CGK9LLR^>
_5E8;&WHB,:\,-Xe8RTZ-Nc<:[<GSL(bR:+>7#@&)#_<Gc#/c60Ce0AX0NSXU(EA
(H<+C[;g2,LW^>87Y>W/TFT4B33M9LDGCf<5?[cR+K71C.0afMBQbf1+]a)K7KT>
0C6U76I\L_I;Z:MR(7cI>B;VMg?d(BfW^HCHZO<&W4\4JQe#02afE(b8U8g^-_W^
/LDEN&A_[=I<#:(J9IO/V=4MC_PHg#0&39W.#\7KdC>1EKV43014H;=_O+C(U<?g
M<KeCXfgCf@D;8bE0TT5RcYG@U]eH?C_2TT),c[.@B@]]bd0BUY0Q/:HA[S:JO.9
GF1SbN6[^CFG1@Nf#VMI._RFZ1Q^X.7,5MW[Ld]G@Ub9G/&LCB70<_AA_NWP(\)N
T-M2eND)T/aNBR?3F:LXQ3A:7f:1c@,I>/[Vde8d()+aCIBRPP[U7+-V+]Z^LH_6
XYUa(Od6UCN^QYdb,C:69P58J0>W^NPOdHZ9)=8aCc(aJ//(/e6Ue/Z]ERIda/2@
G+2,P/Wd2.P3_;;.FT.VJY19I[1S3^316_4VB>@fSaBR]#D82NCU?f5J#;J5g(;I
U2+,PFIH32DT#FU:^/G@DcH=2@(M&dZEbUBaG6\=>bZLJFeK@M;GJ<,bK[6Q>L6M
]4:8b?X/QUb-6ZVZF#+_g?-QG/F3d\4PWZ4R0-O_,W]LFAY9cFA-:H##TaU&cCdB
(V\=M93IU[?7P6;?Q[39SX2,#W<=dG2[+X?GPf&FT96bW#>:Y+F^,/_[DZ9;JDF-
+dT&;f>0&QV2(:2+e@4HBHBgQKH4:VfK,DUS?=-.^8&89d2<_H_IMSGU^(MOO_/;
0&@D4MB,\U.)2D<V2bSZf:UMINM0>[e/bU+c]=(fb5We&1TY(F0S+EO?>>VD[N89
.B:M93DY[;AXK6]QfTEcM[C)HD,\]B>a^)#(5S3B^CV52GE;.dGdO+0?RDT,(Q+G
GS3cc^3V#O,KIX2aP^\fD1e&>S&W^?S.U2<=8:VEH8J>2QIQ^RBS/+8&:d\Q:c<C
ePL4;cZ.,ZZ(O=3D;]H3?3LZ4Q-Y^)Q)G+0HZ5;;f(1PW&]KE;7JcP^YE3MT0fX:
P7),;W@5F@R]PD>]36AE.@3W;7f48gcd1.LL.7V&)-RRf_bX]@)5IY(6_BVFFEJF
IPf3be9.H>MD+7IL+:IXG^?ddCQU1A.Yd.a6=de6e0?W+>O-_aVE4>)+_H)=0fA6
c(?Bb3GU-Zd2X0=E6V?.P9,;O4_G.K43PEF-CIDQAQR:21Fg;SPD?T5UP,d5TB,K
D\6J3A.F(6LdcOe?)IU=GC1==ZQOQA<NdHW&C1&@4#C8g7S58:=[IV=#g/J@5RBN
f@+[B#);JY8&RAdg1DSX^18T)LHE79\1d0E4@>6GFEN-4V&ZL8d[U4G0.>cg>E;A
V(beS9IeT0G./RSfF]QTM8gV8H_d1C1&@:URKW5g_M_#DUFHQ[8R4T^,:905QELR
O[bNW_RbJGQ5XLD]^[6=dV7+@#L(B-9<b58IA.>16Q?Z/KH>=EdF&I8X#7F>V7(D
@?Y^J\V.N//\c21CE#J,_eN#Ed]KG6:Fec#XQ0J2_bLE3@Q.:0)@7g_AL/.-A#AW
75LWBX7GCFE.?I^W<aE(I1)#UQNK<G:#d:Sf+DUX7ag8CI+R5VY:dK,VXBgWS1BK
U0RDI841b&eK7JP:Q.PRgK32e3:0\@@GKc4U/<R]>Tg)5UP+RRBMR.;HVcSC.(T@
<fACOQCW.2G2<B2C+E+S&,D[IHC/?J8S9a1g5HFR?J\?Tf^c6,AN-U8.2?DCOO:6
1\LM.+31fK@9\b7:#K[F5dSZXU9ALJ7#\.NRN6ZdCVN(ef+U+@@<3c?)/>d^_:Gd
=2H?.]\,W6UG?_-P-C;90W-Ce4&LTfC)X;1e)U,WW]Q(1X3gF+(&PR?N#TL:M2[,
#d_)H(ZGE,g\]ME07G(CQXI._AfHLW@S?JGY:81W:_M:_ARBX7JgJ<cH,c)68]d&
Y)2M-4FTYTFUA8E#K1UQI6E=7Ra7S2T=\3O=CS^TdU]_SX/-].;3]b?)Le+0SY?I
=d&+3#P1<G3bZFe1fP((EJDLb2c&:MPJE^(Z)TRS7c\VK9(OT4W#89H4?S?P.K-+
V#0LY7cfa+B.(6\LN2@:M+?gS2IX,D(5RPSGK:>UR0DdZ8WSG66Ub/PL-^F\-7)a
T<Qe,9_AV)&2(Y/[2W?D)CZTJUM&#aA-gaAA:+=GDCfS,GABWS4N\=6S_GY^>Y1Y
8+UW7UIE<,9b[AeL&d<&:dP;GARXCBXe,UOe[\N/EL3eE)Ab)&1Z3ZLU?PWfW#&Z
5_9D6A,0@.;9)=8;8e.EE9WaQH09Q]A<eB;RVGQSM#e0PM_GX5;_5>,=.NKD+.=(
df7?>X7d4?ZTS><+T:EYVBgX>Je@X;F2aZaR64LLQJg<TbG:K23<]5Y#ARDZ@^\;
LNDfdJP7fRT#CUNb##+.,^LPR@OeU^MR#W\@RD?[>YfPfb5(PT[b-B]G[933O)UU
FD+0bSW/HT5L&VR/6b7::V](gP<?GI^Q5BVFWJ(=8]=d#g&/D<FKW8:6[Rf7ZOP8
L\=OGSgdLDO:8fg@-aPa-+]LeM]Rc_KQNV(A(c&1P[73?N=PFgL<X@R\.f,Ug=HR
>^AAP5F2baLd+b_dPOL:-gVa+T.g+fNUWabF-U#9]0JP4AQ9.-^0(AW1cQR,DIV3
W@)>Y(>?7ZT)OLN\UGPf1HXaS@YF_:I&GBg()K+=d-^;NgV=@g]EF/[N/M<&HSc-
/C3@OgB9;D+:cY3>6#/.N.&;/F[6?^B@TFDX/GR-T5EDF4C1([d1?@MBP3CE_9G8
L)eLIPF,Od^K=MKI[[EL/.&/bRFUT#WfQ?Z5f8&5\R&3AYOYTdeUA2a9FKL#7YUV
DW_CYReeZ43B&#YS\CN@M)O?+eD(F@EN0II4g[-F^3_0Rg/C^_Q#eK1gBM?:gO)@
)BC^W2g2IP@+/3L]DU-#?V,O)bD4J#?:g2.9f(15B/9[C/[2DKYRD>b3]?YE,G:0
S98Xd/F9cDbC+AXX17[@)6d>TDCe)AC\]@aGXcg8f-X?,baHD2Y7OW1X9>5XNYbF
D\RUVYDHW4fF8OTGEcC[A:a9:B4dSFUVA(_N)WB4O2O#:X1C]Y+D)1#<8IX_6YNI
MAHDC8e4GT/1O<V./_KDKH6J[6^L1fdYB#OV-P?#FdY74Q>A,/U,5.@ZDdQU0-af
>JCIN\-#@RK#RC?D?\<=]\3aLaJ7FG<7\d@HT3V5cTM@T2()Z4,,Hb]c87UGa3gZ
^#&9#B7(RdFg[I9,3&)V6O]?-=[SID304[H=^F)>TCQZ2^;9S]&,[QOV6(M-8NF[
VO<_K\D\Cc,,]E[3HWL0H/+L6?RL(V;gU2dZgFBQfNI4JB<33.g3SQ):;#0=E#28
b[37XY>A4N(NG6f^PNA.C8(O(R8N2(^/CY0M^<[;JG:Y8<3^#[.5Y.<CDa[[D:#D
L>-f>M1SY7H@]>Y7K5EdI,_M_4g:Wc2XXL;.X:@Qf#ZE0ZE+?[)SE]W52=(PQ[FO
\db-,V5@.:498A.;cZS#\e7^24[Rb7_?7gEO[E)eK\.?dF,ZXW(.^e?\?aF]LH(.
4T<85f3Y#<L8Fa98L3B@Hgb3=b7R?5P\D&VP<J329IJ6YdA&E,Q_3F[Z&3KW,VXC
^:V_b@\LOFb35P=a]6J(Z<^Me)d]#\+OA63NU8.Ha_X.a]P8,[FP7/+YFAL76MEC
5TMA:XM]8g0//>#gSSX_0LIdSbKNb67<=_1]1+MbU-+6,61aQ_J978XMN9/T#5<Q
GYbF4CS90M8=@ZGF77OM7+NcB&HNNcgQ?Qe(g>_/@AMcANF_ZdgY;M^cIADX8[X^
-EF.7Z8G@5AB;R5]2JScfXRDM1Y,91N]d+YgM^\<<+B@)Y?P\ZSFR//+#7]&=4SE
77_Xece,b#,C?2P<2_;U;;+c@91&RL>J)e3B1,NNAGEJ&=?fe>1M;)#572Fea^-b
f\#U?Gbbf74\HDgWB^T?(XH0\O+YDgbD@,F3WZPNZC<Kf#-(,/N0=/BFEQV[SO@3
U@YB=BH20#@J7CT_fZ(>ULXDfZgD#&^TP#T<H3D1AD.9f(;UA8bY=PSV^\,WDMZb
TJ/:gH7+^J8]RE-Ge5-I,,K:#>0.Kfa0JAd49HI><6AfE:3(CB9WU78aU)WgT.UH
/SQF1)RQLS2?>^-74))^&N.XH=;?df-)Ce6V)?1,.6RE8-BgeW(#e.?1=FT:+B+:
[3]-B\bc#N+YO?6DIT.);bZ:.(A<f2=01;S\:U([54fRg;?=<[OF_R5R;^^#/[cK
I0QI2&\J^BJY-IH:cPfJ3(CfOg&,(BFLC5JE1L;JM^AN4=K5F1/_E0,0DRB([g/;
>/JXT8OH.ISV#&gW##A90d&]?^FKB<4T+2XA]a>WN129K6;YYU>;X]A]efT@KO)b
4be#GPL7.W_TaP<5PS3LK]LX4E[S;TJIN6?8^Wb)YW0O#3b#bO4Y@g;46d[bVbe@
+MY,2(;UCMbc9,JW=YR&\\OK9VCfJY^QI)\3KCP3=@Rca^[gE06\Q8&Z8/-]@.S]
1&-W:fbNE[:Y.JNLVFDFZ\Y7Qd?XH.@/6@E^]Y:6^V7Y-AO=^V6=_b.1_6Sb+0CP
Pg_8+,M;Q]X3TWa#TLVHT1#7X::7gP,09PdY?IRH(MBL>Y(8+ZJX8>([F_+UDP/J
]/cg=cA_#E.@fDL>W??J?HVJ0&[@]b)#\C1c03gF8<XC23N@8/R173QJQJe\F@<^
c+]G2#)>f\=e]g>@<eEP9MTR]N8^<aWRWMVCN.Gd8XK4G?#\8gcHUZc0UF+VTA#<
<:XHeKMRK-T09UAYX30#IWXdBDQ.\IE^:2f#.O9CI4Gg@@gBB<QVS<:W3dQcI.dg
_>+S-5,-Y&/6aA;,:JV?]BV1N&9Tb;<GZ^V.Hb\+G&.61b4#92OTVJ@1)a>J(A^?
FAD-Ag@VM63\Yc?@Fe&T\9_eJb+_QS^B\<7QQ99^79-3-c4US-cVDKCY1/Q&JaN#
P-&ZO;1][AfMW_1_6c)C]_/-gJM,LM3Y4e_.@RSGK_-JE8eH-+S?K@SB,5a_3(Q5
?[@dJO3@DR@?T.V@g3U53EI4GT<&g31DXM2Y_C>=P=IDM8QGefTd8GV/N_d<J78X
\CE.f6=f[54(9KD+MU&>W+1]>\Gc]&77>MMg,ISK2]77\]UNYY044:R7d;@T6,Le
f<L>##Z@MPP-H:G>N-<b27c^D9A60P(0D#,7T44JZ;?L;@T>0d<3D3cMX>]]Y^R,
/.CYJDMDD(;C?@8,0^b9C+.d8YA33CX^BK>[6XF\b#2O_UI3,0SPZ(<)JKc9;X9I
4bG@Y1]8F4I1@;#a.=dZ,@Ng(#c88^7.:_d4I?e,&Gb6TdOgbFg<LEeMf2PfC-;T
NM7BUI9:CQ.1Nd6Mf#--@S3R+?B=H9=?H5WK#,+L@_;)gEIAFO5HIa-6:V7UYEPT
\5?(IRZ\HA[\BTU02>&LS^d&bT4W\>Q;aYM3:[1a;C#:;VXTaY=((1ZJ2MP0=E53
K2Z+baJ]UYf7.F&Q3<EY?K-6WR-3N@>+ZZ)aG^NOA+Z#eOURV@30g_R_e--(>fJ,
/M(.L+@-N?O+fB.+K&(dR#Ea/[(V;<IG7J1ZfMMR23<K/F3LS.9A^QASd7(&YTg>
OgRUZbU+E_#a0]VAO/_D+(UD2C^W+S/\0dNfRO^B_ceE@ZN@6.\A6CF70@ST6a]T
JNPID42,fPfd[J@b6/2#.QOYXHOYdY?,Q-&J6V139^TI,@[=LQ3(7GG<UQ&-ZJ:c
^aG^^)Be5Q@<SUKg(LEZ]_IYd;;V[Z3J0Ig4WR>dbQgLcCKR,\]B:J]206bAU1gY
:B=UTOA.9OT.ec,(2:7@+8@-)fgT#Db/4LJP#db3)A5bPTYGQA6O0(&fHb2<SIfc
5L27EX:CGUP3\UdG,MBePBC#H]?C,Y32KZ<L^+CGG8TPfUFH;4fD\A&g9aWK?Z&,
K7e4SA\9O:/Ug8VfB^=GA(M#)E#RHVaNS+PMN;AaU[EF7_\/-9YSa;?P_+EgOg?3
#RHM^RBSJZ,;E0I6;Zb(7D)=40M/9/GNI/A7WRKeULCLXaC2?YC:McLADD_4(ZFa
\00O::BWO6L\+F1)[/[I(5EZgU&.>H>EX=Wb:(LK7f2+JVNcVGB1QE0B&:<K@-).
0IbJIK:LCLKAd:gV\D(4.OJ66O5eC&d-U+K_4VTUU2,_a;F2_OZcK34&9g&]DB@T
C+F5-Q.7a(<SAVd-cc>9\V@;-@?B^Q.gJ.([_HTg@D^\[P)92-LT1:Sf^S,W^>2U
A9a:fQH97c78L6]N)KX4[1H<_fRVDHP(3W5G1&N-[MR67G.:O.GN.4J3=R:B^@B@
9KY0)aY/=Z9HIZ+[@1eVXHg6C)3SG;;]bSgXDaXO/C4Qb0<_]Ia9PONOeJEGQ:G#
FH(&dBZfG0Edb8IBBJ:+QaGAU0FeDXdc7LKERR4.E&#,=N9Wd+9Ea4-WQ_(c>J5?
Q]Sg-K2=\_,6#>I.^>K5BW5OUa<9.>KCJ#/S6EV5VDBEBRV+e=++@ET]\WNTg.W6
H&#T_OU-)STeR0e)6Ze5#VBGgO.AO#&fK<bVI\YM5#L1/9QCL>\2#gR2BQ2=,/RP
9?dI<6F-\WJQ&I&5YU]=e=Ia>d9;5>J,M#9\Q)LV_K=a@EJ2a,><59Ae\B/^)IUD
^@&aGX7W+cb?HXFP?6_G[X:/^)>b+S+I6?#41NH-=bGE&JSJLKcY_c^gZU^#32Se
Y=43B[:1[W[Z,R>2+Nf1bdK[1?0)Z)Y^a.:E7EC@>05I:LdQ@DR?T]T8GP&bXUdB
A&df/1D@\#YJdEd@EeK0D&8]7W3-,6VPO(\@Y1dc9ScS\<AN+3.0Ub3@cf)Oa:f4
f;:8+]7,5&,PQ1RDZ8/9bcA-T-.dZbC[#ZJff^N0^P?O1@:)TZBDK0bQAP9];YFN
C5J9H5>;F;YMWH\0F]Uc_UJZc4)I;IHOKgI669@c:5Z8ICAd@1,8_(@<,]/0UP)&
PKcg:4gL,[:4[6;3O2XfOHV,(@F>OI=D&:g+YcQ75b69(TKK/]T])AM:J[]\0#W?
cLUMcG=;ZAV^f:)c(.7#.6?_M\T2W[F\\XZ(dAgV.QcLC.8fVE<YKE-a,g8INcU?
+3HWfL:b7AQXYV]R_?&@^V7G4RG\N^;_(&5cS(V+_RAXV?6_E/E4<]-SS?0>\MAG
OC\@8[9e_b7F;D&I_JW-O-;077G2-8b_=\L^WdTgRd_I,M[X&_QT-Qa<)8+]Q(JG
,_Eb7gH14U7:_CG?26gc76f?JI<A@67>gNC2:G@[8@gQ[Z0NSU5@Q=:U_+@@gY_g
JV=DOe]&G#P9a+:W.M9<<V>fb]:CYBf94Jd&?0Oa13=:-BKR/AeVPI[0-&)3S;A5
V&ZQU=YY#c#<SdWOU/+AW2^+Fa;f0K]:\5,)A0L:HQ>A:O<#&F9;f0#F.+.IHE>T
E,PFe>Zd\FKNAc4W]C>3&Y^6:-e(Q)FL.(#0e\.B2^R_f8L8:Ce54)+J=,L&4D\Z
N_=.J/Xab_:VA]4@6+RN]T;IRV=XNEf;b0Ge#I3<0N=]>@F^bK^g28Tb#9AgCV._
A/>G4OJS-(==^9W+GgR5#3=IU>WQ:\KfWQKAY]71)Hf\.X-T]H1IXWD?A\<d?^:O
AdaK6BJLW@Q9Xc/TYUDJ?TY5^V=agZRc&:7;84T0G&b-bLKZeMB>V2fN@7@/a<2Y
VbYcP+D.SV8d@,Q\7^OPP&\^fE36gKW2>]Hc,D858<-7.He=]6C=8a;2PSM?Zg#V
CG.RF#I1T\e/6#W)f=NB7-N/6-YZ]d(X,XScMaQ8,TZ1G28)]BW=)Rd21@U?PF]Y
57F@,GaN+^VK)EC=R9VgJ57#EeG58[@SHLX/e6^:e4OUddBFgf3?D_:.0d\B:@7P
A:A52>A5?1>eDP1THbbLBXV>JI)9SZRJJ6HgWHbURQ()GNE-bQLW;2#<Be@adOMO
^#DF6bc8,5ZH9FJ/-)aR(b62@B9O0\3LF&MQeHB&1/248=+VVH9\6]^BN_B]Q@F8
Y.DJ57_[TEV:42;Qb0X6eT8Y:A)7@a&=UB-M3;.##YfQ)#gB+W_\J8LEJPF#8KF-
\CN5RG8g+,e0O<&I521^1>Y?K+GA:@FGc_Ygaa9;/@2H7^)H-)OU4MN@@?,;dDf@
bP/92[^3bM^HOOa\<K7+8]3,eT==-W2bbYG97E&=aPQODM6/L1E80#gH.^3<\g;G
.EE9d)Y79eTW[F.=9O,VD-:L^Sf;M71E[XNF,IeE5XQ.Kc_-M1<L@Ra)?MWK.+f&
c>OWdWe>e\Y,]U<C70a@\0Y[OC;G?EDZb_ONOE=5L?_3#BK[HUR&I-BT5O=1TAFQ
N(]5<95Q(_::9Y2.0.NRK=&b,T9J\-[_,UFb^<LBcHFg1,V,F>D-\V@e2;2X3Pg6
3dTNRMf-2W,56?IQ<930U17M0a:D2I_M^D(\G=UH#+9)EMG0W?Pf]LAH,D,4BY/\
[8f]aUN5@_.BK/RPb\F(>YA)VD=A9c7WL>.:W#>G67MYC]f:L<d<W4B,LNBb[[f]
da==::\d[Eg5NA65GUa7.KI<6G1ZN(B=e35a.cgE?H=?B+.N4bGRaeX8>JeHRbeY
XTPgO8]TE^FV-(DGX66\4g:Rbgbb>0)YPfEec2_ab=c/^6NCS)a\]9Q:Zg75?UgY
4PYA2@PUc3=4P=N=Q?(;c2?@8VG:5IJ:L37ACd3=-C&b#c>HSV][9VP^.)FRL5X2
L,[@ZEV88O5g9A1IY=J0MK5O;/g5E03QFWK;D76dEUT&\Z1B^g#PQ>JYWA^X\3HV
f.;YYP-S(d#6^cQ)HcA.)XH>1RcKaGLgS0<ZK:X<^7O0AJ;(c.<3E-JJ_J]#]U,=
A9_;29:NL#&PVA_ML[0Ya#[VaWYJ\X4KZ<e(0g?NAFCUf\QX)a><3&C7;T]4#K0E
QIRJ]/AW=+_.1fFBRRLe7B<^>PL4OMN&)=D&VbW1>>J??b93.IFNV]AZb6[D6)HW
5ICU:TIb2M.2UKbD&NSWUG@ecQ_YW-ZETO:M@C1TA@)?O1RM2E::NCP.g,3R7S&N
CbJHfGc5SC\AOA&c;R^S4]:::S..]44Sf>?8dK[OS0XLH[W1>Q&[\VfYKOD4<]8S
bb8.,,DX,6/@V&E7_+.I/?OM7WS+T=@H>][DOKXCL1;/^AO54?/YdL7HCWA16TTM
d:,JVgJYW@W@[^_T=a9g/PT-8ZBaa,E<3^1O0M-RE7H)aMa\cQJS>AaV8ZQOUg_U
?SQVE&)ILY+4&C2\+RS]Jd&80J6T9T]<cGP6V].eM0GCf9C1Q^5^FOGN1<755#IG
O5ba1c#ag<9\)D]UT;)\.:EQW,/MS6O_TWH\^agN51.Vf\&6;EN0+5W#>Z)NWP[F
+F>Qg1a2XS@,)7^D)Hc?4^=<2V#_)1.<&)=IVdg-?)[OBdUEe&MZDY=8TGRON-I.
]0#5Y@SO--d10T9OVaTe:777e\a3Ig1MN+e;Zd-9[AUIT&?:@f/>egWW3XI.?NE0
?YUH-e,15_?cNa>bESWZNB(KT-D[46._YU#G7U7&EE0-gf3&I;&Q_#OAAAURd5e7
T4dAZ8W,7PD8O:K788,;S1];FCKT^b6PbN<77<eUJIX&<@Y7cc8]-g?KE=I-6[+e
a;YD<+4?BLJCEXA17JG4?K#P3_KV-E80-LDQa8L6,KOO3/C6B3G4Ng6:\W\IY(]/
9WaM^6b#[2BLc.bKHg7T+XU?>KbXHP3ZgV:9HbU3Q7^4HJE[:]+)e>\V;]=R9H/=
+b@)WVANA?[QQe##&+N.&Q)d(@Ac+43^f>2(<c(/90RVOg<BGQDY.MNUc6,fN[bQ
_9G@=)&Q06#cg-/_d5HZK59232a=Y\MWM,.WH(7.U-T>X.7OcR#2a?bN]Q#;cUP0
-H/A8FgM:A@-.94=\5=ebBSJ?eD:WF:],G&QA,)QH@E3?+C=[Dcdc6SSJJgeHO1J
ABT;IMX3#G^VJ8(J]58Lc3YJ(K4[A7YTD(XYP[c?;&.KC2F#89]4P=.LC\09G4+F
=GV=:8X-^BD]]:4^SNWM3T8eMKT===e+U\#--a3_>ALKP9IbaQ[6U.Q,JK9KOHO0
VN8W/2I#4a2Sf<cRb0_O6/MXRCBUQ1\5F,8-#-_KeC?U.:VfG2(:NQ9eQYTY[I2Z
YVc<7[37WXC:^gR101b5K/4WK4c\&PUa:A#TPS?)9CZ(@ZQ.G20E^g4eO#958VRa
^5:129UI(3=]JIQO8CV,f@4]+89(U)#<W_HQ#FOb<0XfAdQ?Z;FOgQ=CaM:gC8<E
+^+#^:b:@B0\F6)?+A@-6=\[]H@cUbS4<1eGAQDeV3L<=WU9^^bT+Y3e3[LR._;9
177MLCdbW?+8dee9cE@E>E=U?Z&=1)]9\EUb\fQXWAGO0PT31FYWZHM7Xe\]+;;E
D)Q8,0G@555ETZ0:=Rd_M:^L)@a,\4Dd=:LSXPDID3/,L<GI=30EJ&U)^=;^G:Rd
JSG?KZf[9\&@NL&:2:K(6X-W1N83]CPM2=XbONYT9EK-_fZ^cbc2)]\C6b41=VB3
Y+A2f6^_b0[395NaP>O1CMWISE&V3Q1376[=ZPAcWKSV?42?UZae4bVg\bUe\)RG
#6T(/c3bCWeF\7G9?Z5fMRI?[)]C9_BOJ;V7LAFOfRCdF^3\<@JRBeDX2S]3g,-8
N3U)Be4NXB_If]G[(M]W[3G3CA_W:1e8LC043@\Rc##+HSAL/eIQN7W4TeH>_XWg
(S)J[4FCOO<?d=1,Q1+2S+)816:->ZSJ3gd:QaWDg?,G+-^1?B>&:c(B\2DH<=5H
B<_^\?8[>FYSG.CYZI>:4YbCN5<a6?9Le0+<.#,.JdV9Y#G6AB_E2IYb,B_9B7e^
SVCNIe02XS:=;YF\S5OSVeI#ee(+gCJFb4\[:Ub[#bO6U3E,U>5;SC&[YS:(Oab+
UJ17K,MVE7M5^g-@G0VZV/&:NC&L4HX04\=EMf<eXd+-,9LHTP9?#/<S-^0dGb@2
O9-0IS^E:E-<<3]PdU(<+3BG7G3<9T/?ZI8fD-YIfaKW\,2;SK\I-970AA0fG1>>
I8D+0[,eCJ/>\HK]<5:<bQ^QA<,R9JY-:JUa1I\fP#[R+397b9GP@O)21FN@Ed04
K3fZ^YEfX0Ob>IUbbQ<3XBV1_/+P2D\W-Y\2&:D6US=2QM@F.F3g_03+TgcSQF;5
2_:1b^c4/>>D26DV&@((ROG3;M0C9-P0,7MDDJ)T2(5JW?50T>D=SDFBG&SY.L51
7eMHCB4d_f4Va\[RVd,Wb_@;PNf\R4ZNIR(.[:0R^@W;12e\_(X5US24#_7E2K(=
?I)1(8>2EPJW[.-2J]]2Nd^K#XXTbb<QS-d2DP0.0)4W\P8IFG?BfA-++6OA)GSY
#ZOR@Pb^I1;/E]-/^/L5?H\>NS)<(7I@\dQL-&X^9O0[2Q\L-7=Z?7B46LHJNMU&
;\eMLW4P]99-RDdM&NR\XJ#P1;D>W1K-)DAXWVK[Cd1T_dWUHLYV^?S/DVL+7Yg7
b?X(V=2XV,/dXJ\2-Nf^UF0OD.AZbJZ)AB<F42P^I^T0XEI>O.:9\GXd<)@)U/[?
W4&GTFK/fW<eN.[\0d+S\Ce8OLEOM4gQ4Q285-eT66+J&0(gU;+-JZ(2e8NNZ-3>
K;-be@[,NW)[[PaH77TU^(X](JH9631NA9a<+;C#F)/@@#,Ab^Y-:a:NEA+:g,46
DI9(dKPV[OBfMT8HXfC/=O\(V,ZJ?]==FQJJ-#/Z6ecEY:bW0:Z]Y2,eRS/Fc))^
R;Xg)02O_PHGGa^\X:)3#DP(YWLW395XH>]]&c^]4UbF)5\9#<(Tdf)NW2]^Aa4@
BTSc9Zfd<PJd3[\O@B_P=:I6+0dDTD:OKZ-@Ye=JOSE@<]EIMP7-/541&)-Z)NQ@
\3QV;dMR:d,<,FT)R]_RL-?8YS1(@T]Xf\Ef1Z6\7T1=4fI>;R:70+[IR-AJ>Q[8
4?>L@(70F)NP+NKKR;=c+R2LZ9@)DI(&:PD#7+H@^G_5+]__J7:&6C5dIfSA,a#N
Oa+K^)R]]\EIdID3)#G^G]MV/,,>eO6RIK0cP>,IPDQ)_[&OB=5ee(>9cI#[?e91
3\&O1?=YJ[P]d6@(WTC8A&[<M+-gU9YNC52^N7<9S=BB4J5b^UO4K[ag(c1(c:f5
MI]-;/^(AT\YOYcPPME9\/H#S[53BD>b=4Z?#7N/R^TfIY06bZA3gD=F#8)8HNTX
1&dPEE([#RX8#CB6&@81CO-YN1Ffe29\H.T.DBSKHC)B;BL-5+@X7MVKg.X&K>KO
-8M2SP4(/5Y@DV.[.3BMQ?\==<+_;=8KE4&Y5U:eBTN#f@]LS])+gJQV>>5)OU>J
YL/RK4U\KR+0Mb=fO[aWHZVGL_F4?79<Q=c\J@)GEM/_T/6e0ZG])M(c^BRE9cQ^
6;7?:BcJ.ad&(L1()AXbVIb[<cBDg80+G4fT\EV/O/C3WL=&/C5WPQMPf+8Z]8J:
=d_AXN^g6+VO_W;<=cB(;g&>.agC^>H4EN2&a=c;<YReW2gcRa=@._CQX:P?0H/_
0&d,]P))a<U-T7J(I9e@;\@.T;[3J3B55E>74#+1_IV/F>.APd###9\S,[?EN)?g
W0V(cF&2/H#35X+5J7>]5@D@g9\0H(E@d?H97_^:cN?AGHCEKRC<\9a]5Q8+9PQ(
>&H3b1^e?-W<5-bA_ZE.LHcc+R+O&HR7A7:F+X6_dgZ),QJR(=&a9V([O)<;T(ab
D,YLQgPKKQ:d2.KdOg-N--U-,]3[?([\afM[Ib+Baf:LU&19N0_dd(1@3aUXSZV)
K(4Pbb_93>X(R1J]V\&C31_+DMW)>#2,PW:(d:f;BG>EP;@WL=9YK67KD3AOgX+)
X(N,9QWNA5T[B\B]9+fUQ7J_5.:14N:V[A7TZY_(e#IK;P]UY+A:Tb-J-?(ZL61\
UJSPFBYC7-=>J;O,(g[HWH14RNM][//4.]>CIbLBYRWSL0E9.K6WP:ZA6ZT)EG2b
&//O\O/=Ya9HK5Z\XeF1FO<97P]a7C+ca,FZa;/beJ7+U.JJgMS(_[7<:TdP[=53
a^26>3_YP684#2]N?3(-1=7KL1.N<&O)&-YJE)+/9KWRC_B9Wb[BN:fAF+UP.XVb
S@YZT(f:?ZbM\(WBR2-2bP)?=G)M#gW2T1g[/7d12VA><cBf4,Oad:ea?Vg?UZSP
[+HP#&-XWR#B49:e;Q-b(4=#>]1K[<)4085^aTEI^Kda_KNS7e@CKVeUdQac3DYA
<0Z/],JS0>=^J<.GC./=ZSMWEBGWIf-R8B8=++N&^4QZJQZR^Q@+.OBd5-gN\;=J
7#EbXUGV^W1bDDC],))LH6b@0@LX[41dVPVUcScTf,.fLUTdYae-1-N:QXa62?bg
GQVY<CS<,VL04238P78R.@&D;BDMEbT/<2?bGB(?C<=dW;MWZ-9cg/[5+(1dbXTR
4XafI]&[/:K&YM.d&D;WI^HAF?f(b4ST2edc9CE@BC)K\NN3FO@Pc;Ua+FS=;S:E
IUbNAH,D>/ZK.gNMXd3CaNAUO\Ca,a.-f=).)@HCI&JLTUUe5BY,QC6D](MK(4K2
^>00EXf(VHPO&PNfTf<?efGcP\@.U5fc3?egfcf8cRRU,>>U.d6\?AF6gXU=N#H^
OEOG6ZP1Y6?VXd4\0\L?\^1:NRKFVQ?EcLWG\1DR;gD@FaZ,DD+TU([Ne@5Q&]LJ
:UR6Ae[-Bgg7)/Uf67EY@BU;ZTCC.OJ7&PACe;P@9N+MX;SNXURTe;,:bZ2K-1Y8
W.SG\WX/@;#ATYDDaGCc5D4YHB8g6U9WSER08-&RM6S;X&67<V7fWd1K-aPR:SOY
/AL=8G&-b:QMTe[=Q[L&JW+&=7F^d,MP(fT-B[NSX4?.(:6>FM,T_c,UHAQBJ)43
SX:b&TQd[E8eX?=OP\S0<^VdHUO;EJ0MJVMSH6;3(:4,<M.BR##NH[?bbg-1?3.b
S1>3c^_/YbR)YO2M85OEB+O?<5YXE\FU0RY<b[3SBVP&L];<0;f==EgYG0O4Ze,C
E)<RR,GVA@(PS[FGTJ+53799?C7#.PG_O2BJfP6I\U8W&>XG190C&Z@3LEf+P3Y9
ZM?>>-(X1V[fd9#@b?YTB@gYg>N)Q)Z5<#Q7d96X/N?\J\?e21S0DAA(741]Y\_Q
X#Y[.CIf]g+?Sgd.<<M.gNN[3)-bEI\Xg^RWHT/WE&:RQ89,B1<LC6]=eUddPH=d
gQ6C0_B_)M=PLa;+ANO3K2ZI5DO1D2X[I1B&eJ#D0((Odfc+ZUGagXGWTP3gZQJa
Yf3@SZ8JY._>7)\&d4#5^AC&NCK9,BdIGdJ<#)cYXAV_?3YLJ&31[7f#P)UR)C+F
N+:]#Ed0(IZ,J4])BfMg4UbP.K,eF[?O]08>J8a>_U\2;]FBSLL1g:M_(d:AH8^1
ZW-8Bg>SM3)G,R?YJ[9EKe63a:dDJ+#=L+?Q...==7a]<S9?d(f4P^TOHHQ>D<-8
FSd(\g=TC<B6.Qf<CG:#6F8X?I\WZLG5G9@((UMUc.?bKCIY1/RXbV4\e-2R>Wfe
d#\dfa[dC34)F<#86P6<FPeFZf-OM,W3g&WQeDM57H9DFVaa:49dfQ./Y5._+O-V
b/PPAW7:ReSX-7((>;#f754@_QHC30^DedVBI?0<f:Ab#/[-9K5\LZ9K6@-RUgbS
9@YM9GV?Z3CK8e6c8TGCdFSH#9UOR_M:J.JY+3:ERS/@4g=5J8?3LEe_4fF)d;3-
89[I=U.Q9AS>JLI=>:&IN=f<NTS-O2KMDK:B.QS<5@Gb^A/WEN-?5+4fd=-&UPA;
3F-&DPZ]Q<87eMML<HE2bdWFP&QM-<8Y;MAOa154KfL&YZd>b8>F/F/UCU3.\6Va
/6=b[.MZF1V4:eS1+feFOX9M1+0:[M([fg<EV?QA;7]&>YRS\IKL?e/?\.8-,d)_
QC3]8f^&bEBSe/>3/O;&^7Z5_^-)I[)CFAQU#<]HFGIS;44dUH[.OO62:61^5&DG
>YP0U4#[dE\Z]_H&dL/-BY,SFKPPKb@;fe=(>/QA\f(-fda09[YL?)]g]dZI1ONS
)YKDUN/[4?L(7O81R,B6)0NFD1#)DTOVbPFLfcUL/#,]&-C&N9=ZXRcOOQ8<.5c]
WSZW,/g9+><BcL;&JTdfZDM4X7+D2VC)-3S54c).DBR@XIBRSX@X4=:BO1ffJcd(
S]Sb0S;E8R>dg=ELT.4caOD;RX)-c/C._b@3&4Yg&?A#a=:6+N?V9f,\MQG99?B@
]JPZZ\SZ<7@7Ldg)1_(^I=5eKQQMI:E<Ufb0EPZ\EcDKc<&9Q4.M[=9FN/&J.+KS
8)X.cWSf^W+V=O07X9.d495^5,c?gR:3<@b7QcP_C4@bd6_=]YJ<5(JAgOS2U=UL
gb45Z(E^?U3,JJ1>GF0/^gb?1#d[Tg<^@HU]Id4.1ML?]#,U7J<1bNLLONOC5>Tg
0LDceW]<=fcC<-+4Had44HO6aSRBP;3_L.dPS@2(1JA,FR>(X]4AePJSbYQR)d^C
e#+GaN@#>0IO-,(0OJDRY.QfX=aO+[dSEDF<5D8KS+QC+Q=&)=>VG&(B\\OKFRc.
6UAX5<FRb@:2>H6Sb>aAaM)f8U1;4AG@CaB#563D+3,f>P+f4UaZ8NL8SRfYA>@K
g719(R9&683cPB=,X@GC=0KA.5g_^<cegEIe@DJFS;GL5;6=I^UGdS+X51\?K#PM
PLbe^7FS6S_bUZWM07@X20QLE5L&9JJFKL2HCbQ:TAP67PDH/aW52;=MKYRC5[9/
&_W/D_63FNbN22M+32>)JfU?TQ^\-^X8Y>N@XcC@OWU5-\VEM3J?^VR:L)[5aE=S
J6T_DTc9>Vf/8#T+J>,Q/:adaVI6DG@N^NVQdC@YEQaf@LbFB\B4LVaKZJeNXI3a
X23CI(@GYC2?:T]g2Z[G8G[,d&LgV49TCX7gd9IVGON#OY.U#8\F&,e^_JZG<G;9
X^,L=_5_Ze;]<_<@92ANT6^D5g2;>#_70;_FRT&XUM&?GR0W\HKaO,5I&/9UZO(Z
.b>[YVRd/<H3/<+L#Yd3FK?ReYF>ADV[/VC3<PIg#]404d2CD]6A6YRf5IH+HA@F
7Z+/[=^F8R2Q/(U-30+#aJK08(]O;2S9H@SW0+M^#):WVBZK7^D3CU4X\5MJ]>42
FF#-7UJ5CYDBbX_N94g2UM7#I?7Q^;cG+Eb2&M5<GFDSW9XC[1Ef([X:U562D&&7
LM/3NNbJL09ZPSRB>[J[ac.@\E[2L(bC:.^W:2SOSO@(F9<<HF@>YZCU2KVV.(?:
+-GcEI>772ICSB;F60BM,NVcLQL3B=IE<1JTdJ]5X9)#d[_cJce6_WIg78;F_NRf
1F-A_ZfabK36aNR&Bb(O(<[afWM=2/JCA4KA62DU1XQH9WH(d5(8[-QE-I65(SH\
^=D^KSE,^6XC,3\8F[ISJd<R)[(>g?#JFE@QO_;I/,Z_ZW9P(.4_<?0JS-GZCdYH
FJ&c9eVA925KGQgZ@LJS/&a?O(S+:B]-Hf_12,@_CbU2>Z0QFaa,MCLUL\U\96ca
Z=dT]N:U6?aASIb<#P3f86#OXK?Q4Q,F4)=7.B[2E:D>FI)1,_cF>gbUFWD>;_S]
1RRe^@O]JELQJS&;OP-HQ<NVaPD3:&@VFeGMC=+IA0fX\D4.-)Ma_)4A#a;D?=-Y
]\5b_.WBbD#]GFW3<4Wb6]Y7,(21bb\48;-F17dJ.3(V4&\0WH<ZVU,N[Y8]?+;N
_dE2Sa:dEAP&&&+86=6_+EC[2J(M^A@9=_DcH<NYU5LYcU8=^/A4W1d#X?>A6M))
f[+/b+><<C)/e2WN\cDMFPQZD_Q?>?LYG>#0?@T(1-7a&\3/K?QB4A3)Seb(>V3T
H,;2AEMg29Y(3+S=Z<P[Yc,8a(<L#W]PH6JX4OSed\<,9d-:]2dD+99<I-F&)W/P
U7MXUg;Z;CYa]c\M1ZAa4@b227>Y]:QR@.PQ+Gb,M\_73PE>;Vd.2>-\C-Q#YaS^
?VX/>0FA8&5d^C]?3GC=F,8GJ=_AV]K/e_4_)CTM+#V4gUVPAbA\X\7ge)dD3YPg
bJ@G[M-:M@fJ#HM^9Wg9UW3-J>,:=#R-TAN;b,_Cb\O,=O(S+>-9R,\,0)K1Cb]B
TbWHW#5Z63#>CHOZ5[PX:<\N_(=#UPH.f+CQ^WWL,#Q[6L)Ad:MQFXS&^K48GC9^
AbW\ac\Q?@Jg/S_L?C0TUSCD9CYR_M7&0<H]ccG5c^A&\H9BHHGR(9SV_IRSA./R
1dX?e:?M^bRW-JYLg;P_gSb3DX>G\^PIKNHCb78&47)g217@;]VJYX=gR1W[9@G+
cJb:[Q]X;T_\1?f99UB\97@J[fbKK2FM7UVY9ST,.Z.N5QMKKOfV(bPQ0-8fV,W/
Pf(@MWN;.U-c-,CT#J.Oa<>F4.2_JbT4;Fe;:YA_QIF0^[+&cSN0<AEc0YIY=Y-X
EG<AT]-a;#B,ZS_2<a4HI9JgdIV@&d&GQ\6fZe?V.Bbe_d3GM0#KWT/CG_PBD-Lf
3:N_7Yc2HTCHaIAWC;-N/eS4FU#XW6OG20.d=WSV3KL91Z)LAZ522,B.F30DGVJN
EbN):HAWf91GR1S[Hc^b]WOW3XH+4LENa:?#F#X7V&9F6VYNCVHCf9F;<X_W/T8F
T&-5CY>fSMBIR0X/.I.D,-NK:AT@=UgTX,(A1TOEOKd:;4bX]>G(E#MMCR-c_L0W
IZ(F-]OOA8B1(/>.W<CLYd5:E_XJeJ?KKc^&SCg>5.b&Y>\b]I@]4g(NU2N^HJQ&
#AJ&\_5P;5BG45^/0YEKTD,^]VQLK(@?2HN:4bH+b5KB)CJ1If18-198U,/8LXJP
R>93AQ67M1.1JGGJS;+bGD-0OU.^^P_Cd&(?=&3+Dd?3-[T#@K0;Q&DNRD?IW&:.
bMNN9T0cBY.dRHZ-cFP5TNMTgY+a7>LF69#_CDgFgJ8J&;Y4OTBfM-+<K?YOE(f4
D\GB=JP,WQ>36;<P+:Ca1dL9gDNQ=VMH]9NFO5b76<NVdXQWX-<I9Q2P:J1DD^>W
8VR<@-A;Afc)Q>ZJZKadBDE?1)E;D,HbSPH,,VcQ?<L^Y3NR\IYUK40\Z:NKHKBg
g&,d:_V84cbg?+_J2g>@-H.W+.I,^,Vb;[Q,E4&U?^T-35/9&U]@>SDXgbFNCN/\
e?_W_Z=#Q)43T5a0eW/CQ.Ib-];+dUP2O1[OCg?3L2A1Qg7gb/dE]DQR[_V13N?0
1aR1C&]&eI&WLAMdYKf7N<>\#DT7dbFL0BV3#Rd8_0KANH#K(9\(=;KJ=(bNbO;D
AZXcK;\Y<E.079VfaH<E,SGaB8G\dgNZI?aTM\M)bTY3-9BYba/(28C:e(BIDVI5
T2GfC>;aXI:4#=L:3d]-#S_X7+,>:C_^8Z^</@S<HK<NDMCg>LX82WZN\?NB8\W7
Y4Z&>GG849^JQI=42,8X3-Z&QaHVR9;#;V\?[7A(EH[Nd5R=Ce)YZNFZa1TfaZgb
\GQF)bMWUPb\CeV+UgPO:TfU3.KKX(,6cL,;:HT6<,1CaW(5Z,AMKfFAKB^:V_;P
.,SA0?2&--/AaTFL(@G&PSbdO670Y[(c]4gZ81-If8QQEL//VB&#3M@MSM)L]9=;
.Cg8.\7XcJVG_;ZSdESc-FDV^1#ZARg&K.OS[;[XW-V^&\G18E.T^W[JX>(H1^d]
-SZ)<g&),V[b/_[>6XFMQbaQU=/6f#AaOGJWIJZSg_Z1LQXe.gZ\VB(G@3SM_Q]T
@-4T\R(G[RA27:/O41X9BP83?TI:,JTd&?IJC;O=<<.,9.7WX^^g5]R,&5F1T[;.
c(gAJLCNFHK8ZIdQ1QQ+HL,37BJTF/#KA2W9(C];@8+66T3dI.VJS#@9D<Nf9dg5
P1g2S;;_>WHPJME)U5DGD[OFZ-EVR_;Db3P).1ZJ4H)EH^d#ZE[I5KZ&bHF(_]22
UMJ??D0:bMY#d>60,8BZI)^:-Q_@cVXSWPU1\VPAd0UGPPW74:6F#U+cDYKM48>H
;J\/-Ja,eT@<,>D])OKTK>aE1-4.=I(c@@(b,[ffHd81V\g/T87O2=_K\;gE+JR#
4,,NJO(E9H<,Y2&XE?fKQS/9?>KSLOSWR;c(Cf8CKO_d3(Gf;\,7M)agS-eFOZ./
fe4ZQ[C[bG;#Yf5FBSGMe@&)^bBKeQ&Ee#Y-EbYS17?D4/Y,EBO[AZ)af)KdR?Y?
43A=)CcXcM.Y4>.5+eHaMM7_QA5939aG4A&2)Kd>gL]Hb-EbF46UHQ>NBAZ2Og7b
dF_c1_<f+XHe>^3&D8(TD+HbCIS,UPGC^>b)&GVg7&.#0c,\J5AdZ8E/=GJC6O.F
V9D(fLX-^d(K>g1+0g+TD7d(75>:QFcG</T7ZK-+[P51g@R:=OESQQ\ST=DCRA:U
V2P+<M?,,eU:,:W^UR>c=a1.2985/XD=W[0C28/)R5@d_d=PHH?E]fN=NQ[<B?dO
EP[+P>=Rg:gNISET62fR4AZ^\^]B746MY.JTD3Sa/K;@#Ib0-aPe/_EW50#BT1c.
_cK8bMCaM^8d=.EIdLZJ=VNE:/)e;eQbDE^E5>VIKC92cBa>L)K:-?J@&G.(d37.
/bW^g]C\cMgWOCf+e9M&#HCEK<B>D14gLHK,aJ,12DG<\&4<JJAGCCCEeL?KA#/@
_AbZ?O.UB-?0L]@@?>7_/^b2f@G@;#9<;gK=ZeY\@c]Wf>X2T,Z>3beB,b&;b)eC
-aRNTTU^N5-IQBF9#BD)M5bUS.SIJ@C@&=eM@&I[DL.U(=0ZZfO-<4Y-LeWdY&HR
F&cZ57H2dC,EHf=[^=b-;fT+dUeVR<R@D_E4&8CEO#DB1E@P_Fc4-\TDZS3Ld>f+
&1>H^EIC>;0McZ(C[,\)2BCT@a^gCH0^8ceR7Z6R\WOE>6OgH;M:(=3gGRJ61dZF
=[fbU5G\774dbDA)R#C#RXBL#XgSAIT0@]M,<BC5H@MW8bIVc7D#^3N)+0BMY>TM
AZ\@6@P8K,U0]C+QZO:4J?aP?IWG,X<b^CEd@f;1T_(>;;X/K.E#)GU5=ZI.9M?6
[KX&PW5B)].<RI[g?@a4bP99VNCZAV8>+f[+M7TE:/7YE#:WH(FI[P6I&RL)_;[?
__]fbA-ASe40W3Rb\3D>VFW80?F@PV^H^)D/;#d5<D33+3^/TIW#A^T+?:gMW.I:
K#;;DU793cVa+T@@=K:PGF]6U6+Y/0e>[D:4bF:Y+^PX&ddN0&SDAMM)F>P6Gf;a
2NAQNH?f,E)G:GQe@4/@L>S]TE/(Q)dGcWS]Dg8O52XWfg#g-85ZX/eAR=1J__GJ
VDDY.R70=Z&>WD4F@JLSbF[#-S0A=I=4E\+COT62SPS?>C9W#,F(LTI&XdEcGG\X
e(?fO./D55>H[BYQ>TcR_^gV4G[A&8;&VXV[+^PS4Y1F^^+bAQbdT\CW5;4eH>B@
gL8;7aP1T@eHaPZV.CO<[V9#b]a=Y7bI_M:M@gNHW2Y@0E6,.#>H#e\^Ud-/[fWX
\)1CA0MH0(Z/N\TcT6?Hge]-9//IU9b&3KQ@8KRVP44-^adL>-d=B[R4NM=E:ERY
T<@:6ZE);449UW4U[V2a]XUIC8P48)FL)gV<\V@^RcG2MRW:O0aO\RWgY4+@<5.Y
ZXO(X-:CbETK#6]]cX_9F^OG?@[7V=3=7)5:@,B+>XA<V/;R0bT25J7eMJ[?RSYQ
VAB:+d4cL6@ec,_6BIQV1Ga-NY<(G6VPdX,B,<[CJF08\M2?3+aV5[Eg?f/]SX,[
=>D[\aZ:Nb/DA/F^M6Y7[a]T]VeZ8DR;C]CHT^=^-+;/V##B3\d-a6[WS(2a-W:R
OBCI@H)-POFIETGQ013L[]#Jeg0^ICVXgS8LE15;#GYb1OM&SOd8>^WO,NOOTd.;
T#/=X)eM@A:]+:O[UM0@LR\UbSODV@c.?Qc0Q:.UX2@(/+KY7G;/@3EC.+[([.2D
053(,bBG__?18b\,5#51fOM5?b1\TC3;CP&T-fSaI6AcgA+#;T:d=Qba9YIAU9=V
&Kb\6F1Q?BT0>X17?EJLg6c\8[JKPNb5(DcO/R9TFB0[g<Wd:/Bf[+1B:GZNG[:W
@8>LKb&LFaGRCY,SQ?VIM6@LEZ_O6[OREIT9:WC<N>RYG@@,:b@O3Y7SLa>5@FV,
N.+X4_B)W1=WSQf#LZRgX>&Ff6R0Vb]DNYd<X1Cd;9U)e_GXIZ=XXc3J2=d]DD?.
7#7JfD#P]]g\>3K=VD^8?DHD7^cgS>K?TKa2,cT[f]PLdUaVBKB81[9HE3ST^Q&.
3Y]XcK3\NDa.&f].N0@7(E-?6(VSaGT3Q@H^6JZ00]3,R8-Y&ga/e^(#Z=^C2=:/
FGXA5@@1J.=3#7=^fAd+B<6[.3Z5AJaC]+H69CFN+@=P/=?0HWOef[W?-5c),?d]
4+?gc3X\g5A0GHJ,[=b6CXNMObUQ87YQC9G<gXHC]=[_,#7QK)TY(0B#76[gFD)f
4#@V-.-&f[GY[1:0#NQJ9C[A,,U)]?MDVMZCD_a5#0>-,Z<OG&J=CM,HbfG9B][6
Z</1OIb)#B76e?&/KHR3be8YO_8YI;3S6DMC8Y6?AXNUB9K?^(]VILa6&B]O/LX5
fEBH0<\8MTJ.cCC^cWBF]JI(_X^d<[#UB.fa+:be,V\P8cb+6LUN,XH1/ba/W4cY
9f]YT-RHU<E[FWabR(.^ZF[G6WXCW5fKQgB4#BU2f@G.ANeUee\D9bQge=EV=JYE
ed/YK5P5Vb9[KHOAc=_L(_<G];>HTY:^?-71DQ/O(7+&Q.?/>D:.2>RJ6f0QT<U<
7<BU_CcP9=dP04\;[3fg,R]DN?cE#A[8Q2fHF9LB\8_#/]TLB-a8G5A2X_EU\bC(
J5,[g,GD?06ebe;DJKJdW[CVT#^/?3Q[5P?^4,A5D31)3_(R4LB.+fDJ=5d1=:;F
dVND<9EMT+<Q4/?B7Y)S0GbXK9PM@::Y9J:19;_FV]7C[=ec]>=9Y[UJ;&e<PH33
)184P_NdLP#b3Fb71.AZ5aKY)PedJ,URAQZGQ5Z+bXECF$
`endprotected
endmodule

