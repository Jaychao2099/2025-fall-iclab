//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   ICLAB 2025 Fall 
//   Lab11 Exercise : Geometric Transform Engine (GTE)
//   File Name : PATTERN.v
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

`ifdef RTL
    `define CYCLE_TIME  8
    `define GTE_CORE u_GTE
`elsif GATE
    `define CYCLE_TIME  8
    `define GTE_CORE u_GTE
`elsif POST
    `define CYCLE_TIME  20.0
    `define GTE_CORE u_CHIP.CORE
`endif

`define PAT_NUM 10000          // Number of command patterns
`define MAX_LATENCY 5000  // Max latency constraint 

module PATTERN(
    // Output signals
    clk,
    rst_n,
    in_valid_data,
    data,
    in_valid_cmd,
    cmd,    

    // Input signals
    busy
);

// ========================================
// I/O declaration
// ========================================
output reg        clk, rst_n;
output reg        in_valid_data;
output reg  [7:0] data;
output reg        in_valid_cmd;
output reg [17:0] cmd;

input busy;

// ========================================
// clock
// ========================================
real CYCLE = `CYCLE_TIME;
always  #(CYCLE/2.0) clk = ~clk; // Clock generation

// ========================================
// integer & parameter
// ========================================
integer patnum = `PAT_NUM;
integer i_pat;
integer f_in_1, f_out_1;
integer latency;
integer total_latency;
integer i, t;
integer pixel_idx;
integer sram_addr;

// ========================================
// Regs
// ========================================
reg [7:0]   data_temp;
reg [17:0]  cmd_temp;
reg [6:0]   current_md; // Store Destination Index
reg [31:0]  sram_r_data; // Temp storage for wide SRAM data
reg [7:0]   your_ans;
reg [7:0]   golden_ans;

// Dummy register to skip comments in output.txt
reg [8*40:1] str_dummy; 

// ========================================
// Initial Block
// ========================================
initial begin
    // Open input and output files
    // Generated by Python script
    f_in_1  = $fopen("../00_TESTBED/input.txt", "r");
    f_out_1 = $fopen("../00_TESTBED/output.txt", "r");

    if (f_in_1 == 0)    begin $display("Failed to open input.txt");     $finish; end
    if (f_out_1 == 0)   begin $display("Failed to open output.txt");    $finish; end
end

initial begin
    // Initialize signals
    clk = 0;
    rst_n = 1;
    in_valid_data = 0;
    data = 'bx;
    in_valid_cmd = 0;
    cmd = 'bx;
    total_latency = 0;

    // 1. Reset Task
    reset_task;

    // 2. Iterate through patterns
    for (i_pat = 0; i_pat < patnum; i_pat = i_pat + 1) begin
        input_task;
        wait_out_valid_task;
        check_ans_task;
        $display("\033[0;34mPASS PATTERN NO.%4d,\033[m \033[0;32m     Execution Cycle: %3d\033[m", i_pat, latency);
    end

    // 3. Final Pass
    YOU_PASS_task;
end

// ========================================
// Safety Guard
// ========================================
always @(*) begin
    // Busy cannot overlap with input valid signals [cite: 728]
    if ((!busy && in_valid_data) || (!busy && in_valid_cmd)) begin
        $display("----------------------------------------------------------------------------------------------------------------------");
        $display("                                                        FAIL!                                                         ");    
        $display("                                    The busy signal cannot overlap with in_valid.                                     ");
        $display("----------------------------------------------------------------------------------------------------------------------");
        $finish;            
    end    
end

// ========================================
// Tasks
// ========================================

task reset_task; begin 
    rst_n = 1'b1;
    force clk = 0;
    
    // Apply reset
    #CYCLE; rst_n = 1'b0; 
    
    // Reset duration must be 3 times the cycle time 
    #(3.0 * CYCLE);
    
    rst_n = 1'b1;
    
    // Check initial conditions
    // Busy should be reset to 1 after reset is asserted 
    if (busy !== 1'b1) begin
        $display("----------------------------------------------------------------------------------------------------------------------");
        $display("                                                       FAIL!                                                          ");    
        $display("                                busy signals should be 1 after initial RESET at %8t ", $time);
        $display("----------------------------------------------------------------------------------------------------------------------");
        $finish;
    end
    
    #CYCLE; release clk;
end endtask

task input_task; begin
    // ==========================================
    // Phase 1: Load Image Data (Only at Start)
    // ==========================================
    // "in_valid_data will come after reset" [cite: 715]
    if (i_pat == 0) begin
        @(negedge clk); 
        $display("Loading 128 Images into GTE...");
        
        in_valid_data = 1'b1;
        // 128 images * 16 * 16 = 32768 cycles continuously [cite: 716]
        for (i = 0; i < 32768; i = i + 1) begin
            t = $fscanf(f_in_1, "%h", data_temp); 
            data = data_temp;
            @(negedge clk);
        end
        in_valid_data = 1'b0;
        data = 'bx;
        $display("Image Loading Complete.");
    end

    // ==========================================
    // Phase 2: Send Command
    // ==========================================
    // "The first command will come in 2~4 negative edge of clock after in_valid_data falls" 
    // "The next command will come in 2~4 negative edge of clock after busy falls" 
    
    t = $urandom_range(2, 4);
    repeat (t) @(negedge clk);

    // Read Command
    t = $fscanf(f_in_1, "%h", cmd_temp);
    
    // Store Destination Index for checking answer later
    // Format: {opcode(2), funct(2), ms(7), md(7)}
    current_md = cmd_temp[6:0]; 

    in_valid_cmd = 1'b1;
    cmd = cmd_temp;
    @(negedge clk); // Delivered for only one cycle [cite: 721]
    
    in_valid_cmd = 1'b0;
    cmd = 'bx;
end endtask

task wait_out_valid_task; begin
    latency = 0;
    // Latency is clock cycles between falling edge of in_valid_cmd and negative edge of busy falling 
    while (busy !== 1'b0) begin
        latency = latency + 1;
        if (latency > `MAX_LATENCY) begin
            $display("----------------------------------------------------------------------------------------------------------------------");
            $display("                                                       FAIL!                                                          ");
            $display("                                    The execution latency exceeded %d cycles                                          ", `MAX_LATENCY);
            $display("----------------------------------------------------------------------------------------------------------------------");
            $finish;
        end
        @(negedge clk);
    end
    total_latency = total_latency + latency;
end endtask

task check_ans_task; begin
    // Skip comment line in output.txt if present (e.g., "// Cmd 0: MX...")
    // Adjust logic if your Python script output format differs
    // Assuming format: // Cmd N: OP Src=X Dst=Y
    t = $fscanf(f_out_1, "%s", str_dummy); 
    // $display("str_dummy=%s, i_pat=%d, current_md=%d", str_dummy, i_pat, current_md);
    // Consume the rest of the line until newline if needed, depends on file content
    // Here we assume fscanf reads string by string. We read 5 strings to skip header.
    t = $fscanf(f_out_1, "%s", str_dummy);
    t = $fscanf(f_out_1, "%s", str_dummy);
    // $display("t=%s, i_pat=%d, current_md=%d", str_dummy, i_pat, current_md);
    t = $fscanf(f_out_1, "%s", str_dummy);
    // $display("t=%s, i_pat=%d, current_md=%d", str_dummy, i_pat, current_md);
    t = $fscanf(f_out_1, "%s", str_dummy);
    // $display("t=%s, i_pat=%d, current_md=%d", str_dummy, i_pat, current_md);
    t = $fscanf(f_out_1, "%s", str_dummy);
    // $display("t=%s, i_pat=%d, current_md=%d", str_dummy, i_pat, current_md);

    // "Pattern will only fetch the image[md] stored in SRAM and check answer" [cite: 672]
    // "TA will check the values of destination images stored in SRAM when your busy is low" [cite: 677]
    for (pixel_idx = 0; pixel_idx < 256; pixel_idx = pixel_idx + 1) begin
        
        // Read Golden Answer
        t = $fscanf(f_out_1, "%d", golden_ans);
        // $display("golden_ans=%d, i_pat=%d, current_md=%d, pixel_idx=%d", golden_ans, i_pat, current_md, pixel_idx);

        // Fetch Your Answer from SRAM (Backdoor Access)
        // Adjust hierarchy path (u_GTE) if necessary
        
        if (current_md < 16) begin 
            // MEM0 (Img 0-15) - 8-bit
            sram_addr = current_md * 256 + pixel_idx;
            your_ans = `GTE_CORE.MEM0.Memory[sram_addr]; 
        end 
        else if (current_md < 32) begin
            // MEM1 (Img 16-31) - 8-bit
            sram_addr = (current_md - 16) * 256 + pixel_idx;
            your_ans = `GTE_CORE.MEM1.Memory[sram_addr];
        end
        else if (current_md < 48) begin
            // MEM2 (Img 32-47) - 8-bit
            sram_addr = (current_md - 32) * 256 + pixel_idx;
            your_ans = `GTE_CORE.MEM2.Memory[sram_addr];
        end
        else if (current_md < 64) begin
            // MEM3 (Img 48-63) - 8-bit
            sram_addr = (current_md - 48) * 256 + pixel_idx;
            your_ans = `GTE_CORE.MEM3.Memory[sram_addr];
        end
        else if (current_md < 80) begin
            // MEM4 (Img 64-79) - 16-bit
            // Addr 0 -> {pixel0, pixel1} (Big Endian per Fig 19) [cite: 631]
            sram_addr = (current_md - 64) * 128 + (pixel_idx / 2);
            sram_r_data = `GTE_CORE.MEM4.Memory[sram_addr]; 
            
            if (pixel_idx % 2 == 0) your_ans = sram_r_data[15:8];
            else                    your_ans = sram_r_data[7:0];
        end
        else if (current_md < 96) begin
            // MEM5 (Img 80-95) - 16-bit
            sram_addr = (current_md - 80) * 128 + (pixel_idx / 2);
            sram_r_data = `GTE_CORE.MEM5.Memory[sram_addr];
            
            if (pixel_idx % 2 == 0) your_ans = sram_r_data[15:8];
            else                    your_ans = sram_r_data[7:0];
        end
        else if (current_md < 112) begin
            // MEM6 (Img 96-111) - 32-bit
            // Addr 0 -> {p0, p1, p2, p3} (Big Endian per Fig 20) [cite: 652]
            sram_addr = (current_md - 96) * 64 + (pixel_idx / 4);
            sram_r_data = `GTE_CORE.MEM6.Memory[sram_addr]; 
            
            case (pixel_idx % 4)
                0: your_ans = sram_r_data[31:24];
                1: your_ans = sram_r_data[23:16];
                2: your_ans = sram_r_data[15:8];
                3: your_ans = sram_r_data[7:0];
            endcase
        end
        else begin
            // MEM7 (Img 112-127) - 32-bit
            sram_addr = (current_md - 112) * 64 + (pixel_idx / 4);
            sram_r_data = `GTE_CORE.MEM7.Memory[sram_addr];
            
            case (pixel_idx % 4)
                0: your_ans = sram_r_data[31:24];
                1: your_ans = sram_r_data[23:16];
                2: your_ans = sram_r_data[15:8];
                3: your_ans = sram_r_data[7:0];
            endcase
        end

        // Compare
        if (golden_ans !== your_ans) begin
            $display("************************************************************"); 
            $display("                    FAIL at Pattern %d                      ", i_pat);
            $display(" Destination Index (md): %d", current_md);
            $display(" Pixel Coordinate: (%2d, %2d) (Index: %3d)", pixel_idx/16, pixel_idx%16, pixel_idx);
            $display(" SRAM Address: %d", sram_addr);
            $display(" Expected: %3d (Hex: %2h)", golden_ans, golden_ans);
            $display(" Received: %3d (Hex: %2h)", your_ans, your_ans);
            $display("************************************************************");
            repeat (2) @(negedge clk);
            $finish;
        end
    end
end endtask

task YOU_PASS_task; begin
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                  Congratulations!                                                    ");
    $display("                                           You have passed all patterns!                                              ");
    $display("                                           Total Latency = %d cycles", total_latency);
    $display("                                           Clock Period  = %.1f ns", CYCLE);
    $display("                                           Total Time    = %.1f ns", total_latency * CYCLE);
    // Performance = Chip area * Total latency 
    // Note: Area is calculated after synthesis, so only Latency is shown here.
    $display("----------------------------------------------------------------------------------------------------------------------");
    repeat (2) @(negedge clk);
    $finish;
end endtask

endmodule



// //++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
// //   ICLAB 2025 Fall 
// // Lab11 Exercise : Geometric Transform Engine (GTE)
// //      File Name : GTE.v
// //    Module Name : GTE
// //++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

// `ifdef RTL
// 	`define CYCLE_TIME  20.0
// `elsif GATE
//     `define CYCLE_TIME  20.0
// `elsif POST
//     `define CYCLE_TIME  20.0
// `endif

// // `define PAT_NUM 99      // Number of patterns
// `define MAX_LATENCY 100 // Max latency for each pattern
// // `define OUT_NUM 3       // The number of output for each pattern

// module PATTERN(
//     // Output signals
//     clk,
//     rst_n,
	
//     in_valid_data,
// 	data,
	
//     in_valid_cmd,
//     cmd,    

//     // Input signals
// 	busy
// );

// // ========================================
// // I/O declaration
// // ========================================
// // Output
// output reg        clk, rst_n;
// output reg        in_valid_data;
// output reg  [7:0] data;
// output reg        in_valid_cmd;
// output reg [17:0] cmd;

// // Input
// input busy;

// // ========================================
// // clock
// // ========================================
// real CYCLE = `CYCLE_TIME;
// always	#(CYCLE/2.0) clk = ~clk; //clock

// // ========================================
// // integer & parameter
// // ========================================
// integer patnum = `PAT_NUM;
// integer i_pat, a;
// integer f_in_1, f_in_2;
// integer f_out_1, f_out_2;
// integer latency;
// integer total_latency;
// integer i;
// integer out_num;

// // ========================================
// // wire & reg
// // ========================================
// // reg  []  in_1_reg;
// // reg  []  in_2_reg;
// reg  [7:0]  golden_out_1[0:255];
// // reg  []  golden_out_2;

// //================================================================
// // design
// //================================================================

// /*
// You should fetch the data in SRAMs first and then check answer!
// Example code:
// 	golden_ans = u_GTE.MEM7.Memory[ 5 ];  (used in 01_RTL / 03_GATE simulation)
// 	golden_ans = u_CHIP.MEM7.Memory[ 5 ]; (used in 06_POST simulation)
// */

// initial begin
//     // Open input and output files
//     f_in_1  = $fopen("../00_TESTBED/input.txt", "r");
//     f_out_1 = $fopen("../00_TESTBED/output.txt", "r");
//     // f_in_2  = $fopen("../00_TESTBED/input2.txt", "r");
//     // f_out_2 = $fopen("../00_TESTBED/output2.txt", "r");

//     if (f_in_1 == 0)    begin $display("Failed to open in_1_file.txt");     $finish; end
//     if (f_out_1 == 0)   begin $display("Failed to open out_1_file.txt");    $finish; end
//     // if (f_in_2 == 0)    begin $display("Failed to open in_2_file.txt");     $finish; end
//     // if (f_out_2 == 0)   begin $display("Failed to open out_2_file.txt");    $finish; end
// end


// initial begin
//     // Initialize signals
//     reset_task;

//     // Iterate through each pattern
//     for (i_pat = 0; i_pat < patnum; i_pat = i_pat + 1) begin
//         input_task;
//         wait_out_valid_task;
//         check_ans_task;
//         $display("\033[0;34mPASS PATTERN NO.%4d,\033[m \033[0;32m     Execution Cycle: %3d\033[m", i_pat, latency);
//     end

//     // All patterns passed
//     YOU_PASS_task;
// end



// always @(*) begin
//     if ((busy && in_valid_data) || (busy && in_valid_cmd)) begin
//         $display("----------------------------------------------------------------------------------------------------------------------");
//         $display("                                                        FAIL!                                                       ");    
//         $display("                                    The busy signal cannot overlap with in_valid.                                     ");
//         $display("----------------------------------------------------------------------------------------------------------------------");
//         $finish;            
//     end    
// end

// task reset_task; 
// begin 
//     rst_n           = 1'b1;
//     in_valid        = 1'b0;
//     total_latency   = 0;
//     // golden_out_1    = 0;
//     // golden_out_2    = 0;
//     integer m;
//     for (m = 0; m < 256; m = m + 1) begin
//         golden_out_1[m] = 0;
//     end

//     force clk = 0;

//     // Apply reset
//     #CYCLE; rst_n = 1'b0; 
//     #CYCLE; rst_n = 1'b1;
//     // Check initial conditions
//     if (busy !== 'd1) begin
//         $display("----------------------------------------------------------------------------------------------------------------------");
//         $display("                                                       FAIL!                           ");    
//         $display("                               busy signals should be 1 after initial RESET at %8t ", $time);
//         $display("----------------------------------------------------------------------------------------------------------------------");
//         repeat (2) #CYCLE;
//         $finish;
//     end
//     #CYCLE; release clk;
// end 
// endtask

// task input_task; begin
//     // repeat (5) @(negedge clk);
//     // a = $fscanf(f_in, "%s", in_1);
//     // a = $fscanf(f_in, "%s", in_2);
        
//     // in_valid = 1'b1;
//     // for(i = 0 ; i <  ; i = i + 1) begin
//     //     a = $fscanf(f_in_1, "%h", in_1_reg);
//     //     a = $fscanf(f_in_2, "%h", in_2_reg);

//     //     in_1 = in_1_reg;
//     //     in_2 = in_2_reg;
        
//     //     @(negedge clk);
//     //     in_1    = 'bx;
//     //     in_2    = 'bx;
//     // end
//     // in_valid = 1'b0;
// end endtask

// task wait_out_valid_task; begin
//     latency = 0;
//     while (busy !== 1'b0) begin
//         latency = latency + 1;
//         if (latency == `MAX_LATENCY) begin
//             $display("----------------------------------------------------------------------------------------------------------------------");
//             $display("                                                    FAIL!                           ");
//             $display("                            The execution latency exceeded %d cycles at %8t   ", `MAX_LATENCY, $time);
//             $display("----------------------------------------------------------------------------------------------------------------------");
//             repeat (2) @(negedge clk);
//             $finish;
//         end
//         @(negedge clk);
//     end
//     total_latency = total_latency + latency;
// end endtask

// task check_ans_task; begin
//     // Initialize output count
//     // out_num = 0;
    
//     a = $fscanf(f_out_1, "%s", golden_result1);
//     // a = $fscanf(f_out_2, "%s", golden_result2);
    
//     // Only perform checks when out_valid is high
//     while (out_valid === 1) begin
//         a = $fscanf(f_out_1, "%s", golden_result1);
//         // a = $fscanf(f_out_2, "%s", golden_result2);

//         // Compare expected and received values
//         if (out_1 !== golden_result1) begin
//             $display("************************************************************");  
//             $display("                          FAIL!                           ");
//             $display(" Expected:  = %d, = %d", golden_result1, golden_result2);
//             $display(" Received:  = %d, = %d", out_1, out_2);
//             $display("************************************************************");
//             repeat (9) @(negedge clk);
//             $finish;
//         end else begin
//             @(negedge clk);
//             // out_num = out_num + 1;
//         end
//     end

//     // // Check if the number of outputs matches the expected count
//     // if(out_num !== `OUT_NUM) begin
//     //     $display("************************************************************");  
//     //     $display("                          FAIL!                              ");
//     //     $display(" Expected one valid output, but found %d", out_num);
//     //     $display("************************************************************");
//     //     repeat(9) @(negedge clk);
//     //     $finish;
//     // end
// end endtask

// task YOU_PASS_task; begin
//     $display("----------------------------------------------------------------------------------------------------------------------");
//     $display("                                                  Congratulations!                                                    ");
//     $display("                                           You have passed all patterns!                                               ");
//     $display("                                           Your execution cycles = %5d cycles                                          ", total_latency);
//     $display("                                           Your clock period = %.1f ns                                                 ", CYCLE);
//     $display("                                           Total Latency = %.1f ns                                                    ", total_latency * CYCLE);
//     $display("----------------------------------------------------------------------------------------------------------------------");
//     repeat (2) @(negedge clk);
//     $finish;
// end endtask

// endmodule



